#Software: 1.4.5-unstable-66-4e44b43 (commit 4e44b43)
#Command: /home/cuser/programs/breakdancer/breakdancer-max -q 10 D00-123546_S1_L001_.breakdancer_config.txt 
#Library Statistics:
#D00-123546_S1_L001_.bwa.drm.sorted.bam	mean:160	std:50	uppercutoff:310	lowercutoff:10	readlen:150	library:D00-123546_S1_L001_	reflen:0	seqcov:0	phycov:-nan
#Chr1	Pos1	Orientation1	Chr2	Pos2	Orientation2	Type	Size	Score	num_Reads	num_Reads_lib	D00-123546_S1_L001_.bwa.drm.sorted.bam
