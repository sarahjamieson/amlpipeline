#Software: 1.4.5-unstable-66-4e44b43 (commit 4e44b43)
#Command: /home/cuser/programs/breakdancer/breakdancer-max -q 10 04-.breakdancer_config.txt 
#Library Statistics:
#04-.bwa.drm.sorted.bam	mean:160	std:50	uppercutoff:310	lowercutoff:10	readlen:150	library:04-	reflen:3015834171	seqcov:0.0193844	phycov:0.0103383	1:4	2:49252	4:13481	8:10	32:42
#Chr1	Pos1	Orientation1	Chr2	Pos2	Orientation2	Type	Size	Score	num_Reads	num_Reads_lib	04-.bwa.drm.sorted.bam
chr1	11073698	4+0-	chr1	11073793	6+7-	DEL	210	99	4	04-.bwa.drm.sorted.bam|4	2769.46
chr1	27533863	2+0-	chr1	27533919	87+86-	DEL	215	99	85	04-.bwa.drm.sorted.bam|85	276.36
chr1	27534964	9+5-	chr1	27535008	9+5-	DEL	159	99	3	04-.bwa.drm.sorted.bam|3	NA
chr1	27535153	9+5-	chr1	27535155	0+3-	DEL	186	99	3	04-.bwa.drm.sorted.bam|3	1052.81
chr1	33670863	2+0-	chr1	33670879	0+2-	DEL	183	97	2	04-.bwa.drm.sorted.bam|2	192.25
chr1	36931415	4+0-	chr1	36932128	37+25-	ITX	-11	99	13	04-.bwa.drm.sorted.bam|13	390.71
chr1	36931983	37+25-	chr1	36932038	0+4-	DEL	195	99	4	04-.bwa.drm.sorted.bam|4	3658.05
chr1	36932128	37+25-	chr1	36932144	67+36-	DEL	181	99	21	04-.bwa.drm.sorted.bam|21	6921.11
chr1	36933183	67+36-	chr1	36933236	8+9-	DEL	176	99	6	04-.bwa.drm.sorted.bam|6	23652.57
chr1	43814823	4+3-	chr1	43814889	4+3-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	NA
chr1	43814942	6+4-	chr1	43815095	6+4-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr1	115256219	15+0-	chr1	115256271	15+18-	DEL	194	99	14	04-.bwa.drm.sorted.bam|14	16666.86
chr1	115256467	15+18-	chr1	115256554	1+5-	DEL	228	99	4	04-.bwa.drm.sorted.bam|4	4803.01
chr1	115256612	15+18-	chr1	115256722	0+2-	DEL	285	81	2	04-.bwa.drm.sorted.bam|2	3034.58
chr1	115258468	39+30-	chr1	115259001	39+30-	DEL	200	99	24	04-.bwa.drm.sorted.bam|24	NA
chr1	188869503	5+0-	chr1	188870048	18+15-	ITX	-11	99	7	04-.bwa.drm.sorted.bam|7	993.90
chr1	188869695	3+0-	chr1	188869763	18+15-	DEL	162	99	3	04-.bwa.drm.sorted.bam|3	6600.22
chr1	188869903	18+15-	chr1	188869986	0+3-	DEL	173	99	3	04-.bwa.drm.sorted.bam|3	1491.70
chr1	188870048	18+15-	chr1	188870072	0+3-	DEL	231	99	3	04-.bwa.drm.sorted.bam|3	1007.34
chr2	4561398	4+0-	chr2	4561522	44+43-	DEL	222	99	38	04-.bwa.drm.sorted.bam|38	374.43
chr2	4561955	44+43-	chr2	4562049	0+2-	DEL	275	72	2	04-.bwa.drm.sorted.bam|2	164.64
chr2	25456956	4+0-	chr2	25457002	3+6-	DEL	224	99	4	04-.bwa.drm.sorted.bam|4	4456.55
chr2	25456902	3+0-	chr2	25457002	3+6-	DEL	165	92	2	04-.bwa.drm.sorted.bam|2	7273.89
chr2	25457205	7+5-	chr2	25457363	7+5-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	NA
chr2	25458489	5+0-	chr2	25458503	6+9-	DEL	207	99	5	04-.bwa.drm.sorted.bam|5	3017.41
chr2	25459822	8+4-	chr2	25460032	8+4-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	25461700	2+0-	chr2	25462165	6+5-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	599.09
chr2	25462165	6+5-	chr2	25462172	1+2-	DEL	187	88	2	04-.bwa.drm.sorted.bam|2	7534.55
chr2	25462071	2+2-	chr2	25462083	2+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	25463091	41+26-	chr2	25463763	41+26-	ITX	-13	99	12	04-.bwa.drm.sorted.bam|12	NA
chr2	25466560	3+0-	chr2	25466604	1+3-	DEL	203	99	3	04-.bwa.drm.sorted.bam|3	1719.60
chr2	25466683	6+4-	chr2	25466744	6+4-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr2	25468260	6+2-	chr2	25468272	1+3-	DEL	184	99	3	04-.bwa.drm.sorted.bam|3	6604.57
chr2	25468849	7+1-	chr2	25469394	8+5-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	1590.23
chr2	25469360	21+10-	chr2	25469788	21+10-	ITX	-12	99	6	04-.bwa.drm.sorted.bam|6	NA
chr2	25470742	11+4-	chr2	25470837	11+4-	ITX	-13	99	3	04-.bwa.drm.sorted.bam|3	NA
chr2	25470837	11+4-	chr2	25470952	35+25-	DEL	202	99	18	04-.bwa.drm.sorted.bam|18	7805.47
chr2	25471408	35+25-	chr2	25471504	0+3-	DEL	217	98	3	04-.bwa.drm.sorted.bam|3	483.64
chr2	25472575	16+8-	chr2	25472689	16+8-	DEL	178	99	5	04-.bwa.drm.sorted.bam|5	NA
chr2	25474918	3+0-	chr2	25474960	0+4-	DEL	188	99	3	04-.bwa.drm.sorted.bam|3	1655.23
chr2	25498276	5+2-	chr2	25498336	5+2-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	25505131	4+0-	chr2	25505148	4+4-	DEL	175	99	3	04-.bwa.drm.sorted.bam|3	1241.93
chr2	25505451	14+3-	chr2	25505612	14+3-	ITX	-15	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	25505612	14+3-	chr2	25505689	0+5-	DEL	177	99	5	04-.bwa.drm.sorted.bam|5	4421.82
chr2	67047071	9+0-	chr2	67047216	5+12-	DEL	180	99	8	04-.bwa.drm.sorted.bam|8	3202.01
chr2	67047155	3+0-	chr2	67047216	5+12-	DEL	166	99	3	04-.bwa.drm.sorted.bam|3	3044.53
chr2	67047645	2+3-	chr2	67047674	2+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	67049333	5+2-	chr2	67049427	5+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr2	99718314	72+53-	chr2	99718880	72+53-	DEL	208	99	51	04-.bwa.drm.sorted.bam|51	NA
chr2	99718880	72+53-	chr2	99718941	10+9-	DEL	204	99	7	04-.bwa.drm.sorted.bam|7	3044.53
chr2	99719068	10+9-	chr2	99719194	0+4-	DEL	182	99	3	04-.bwa.drm.sorted.bam|3	4544.65
chr2	172533772	2+0-	chr2	172533820	0+2-	DEL	205	99	2	04-.bwa.drm.sorted.bam|2	641.51
chr2	198244271	63+53-	chr2	198244659	63+53-	DEL	229	99	47	04-.bwa.drm.sorted.bam|47	NA
chr2	198266124	168+129-	chr2	198267082	168+129-	DEL	218	99	126	04-.bwa.drm.sorted.bam|126	NA
chr2	198267082	168+129-	chr2	198267190	138+114-	DEL	226	99	100	04-.bwa.drm.sorted.bam|100	10747.48
chr2	198267928	138+114-	chr2	198268003	0+5-	DEL	284	99	5	04-.bwa.drm.sorted.bam|5	412.70
chr2	204637047	2+0-	chr2	204637080	59+21-	DEL	191	99	18	04-.bwa.drm.sorted.bam|18	173.89
chr2	204637370	59+21-	chr2	204637428	0+33-	DEL	241	99	33	04-.bwa.drm.sorted.bam|33	2401.51
chr2	209112824	6+0-	chr2	209112924	88+65-	DEL	219	99	56	04-.bwa.drm.sorted.bam|56	1702.40
chr2	209113592	88+65-	chr2	209113702	0+2-	DEL	242	66	2	04-.bwa.drm.sorted.bam|2	281.39
chr2	239140530	6+5-	chr2	239140605	6+5-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr2	239140605	6+5-	chr2	239140718	0+2-	DEL	168	89	2	04-.bwa.drm.sorted.bam|2	3150.06
chr3	983221	2+0-	chr3	983350	4+2-	DEL	205	88	2	04-.bwa.drm.sorted.bam|2	359.92
chr3	32160184	4+0-	chr3	32160198	0+3-	DEL	178	99	3	04-.bwa.drm.sorted.bam|3	486.68
chr3	38181932	4+1-	chr3	38182000	30+11-	DEL	176	99	7	04-.bwa.drm.sorted.bam|7	25648.63
chr3	38182000	30+11-	chr3	38182811	23+11-	ITX	-11	99	7	04-.bwa.drm.sorted.bam|7	286.25
chr3	38182403	23+11-	chr3	38183016	16+7-	ITX	-11	99	5	04-.bwa.drm.sorted.bam|5	1009.88
chr3	56467300	3+0-	chr3	56467333	0+3-	DEL	194	99	3	04-.bwa.drm.sorted.bam|3	86.95
chr3	89905544	20+0-	chr3	89905596	13+33-	DEL	204	99	31	04-.bwa.drm.sorted.bam|31	9523.92
chr3	105438895	117+94-	chr3	105439533	117+94-	DEL	215	99	81	04-.bwa.drm.sorted.bam|81	NA
chr3	105452533	2+0-	chr3	105452589	76+76-	DEL	216	99	71	04-.bwa.drm.sorted.bam|71	1105.46
chr3	106823929	14+8-	chr3	106824134	14+8-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr3	106825397	19+8-	chr3	106825593	19+8-	DEL	177	99	6	04-.bwa.drm.sorted.bam|6	NA
chr3	106825593	19+8-	chr3	106825645	2+7-	DEL	190	99	7	04-.bwa.drm.sorted.bam|7	18452.60
chr3	106825738	19+8-	chr3	106825809	0+2-	DEL	228	75	2	04-.bwa.drm.sorted.bam|2	10819.13
chr3	128199943	20+4-	chr3	128200068	20+4-	ITX	-13	99	4	04-.bwa.drm.sorted.bam|4	NA
chr3	128200213	20+4-	chr3	128200214	1+10-	DEL	171	99	10	04-.bwa.drm.sorted.bam|10	10918.26
chr3	128200650	9+4-	chr3	128200708	9+4-	ITX	-13	99	3	04-.bwa.drm.sorted.bam|3	NA
chr3	128202470	4+0-	chr3	128202563	7+9-	DEL	168	99	6	04-.bwa.drm.sorted.bam|6	6490.09
chr3	128204597	6+1-	chr3	128204683	8+7-	DEL	170	99	4	04-.bwa.drm.sorted.bam|4	10077.64
chr3	128204939	2+3-	chr3	128204954	2+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr3	128205091	18+7-	chr3	128205357	18+7-	ITX	-14	99	5	04-.bwa.drm.sorted.bam|5	NA
chr3	128205357	18+7-	chr3	128205409	37+19-	DEL	195	99	12	04-.bwa.drm.sorted.bam|12	2678.60
chr3	128205915	37+19-	chr3	128205978	2+14-	DEL	204	99	13	04-.bwa.drm.sorted.bam|13	15476.37
chr3	147308554	9+0-	chr3	147308621	20+12-	DEL	195	99	7	04-.bwa.drm.sorted.bam|7	2078.92
chr3	147308699	9+0-	chr3	147308910	0+17-	DEL	329	83	2	04-.bwa.drm.sorted.bam|2	7433.88
chr3	147308792	20+12-	chr3	147308910	0+17-	DEL	213	99	15	04-.bwa.drm.sorted.bam|15	1705.02
chr3	149656432	6+0-	chr3	149656532	42+17-	DEL	219	99	13	04-.bwa.drm.sorted.bam|13	1083.35
chr3	149656755	42+17-	chr3	149656816	0+27-	DEL	243	99	26	04-.bwa.drm.sorted.bam|26	2790.82
chr3	164745395	2+0-	chr3	164745418	2+2-	DEL	186	97	2	04-.bwa.drm.sorted.bam|2	736.97
chr4	55140761	3+0-	chr4	55140862	80+72-	DEL	220	99	64	04-.bwa.drm.sorted.bam|64	919.39
chr4	55143618	2+0-	chr4	55143747	47+32-	DEL	223	99	28	04-.bwa.drm.sorted.bam|28	119.97
chr4	55144332	47+32-	chr4	55144358	0+6-	DEL	238	99	6	04-.bwa.drm.sorted.bam|6	1719.60
chr4	55151917	3+0-	chr4	55151938	20+3-	DEL	195	91	2	04-.bwa.drm.sorted.bam|2	3356.32
chr4	55152029	20+3-	chr4	55152105	9+8-	DEL	197	99	7	04-.bwa.drm.sorted.bam|7	9367.28
chr4	55152377	9+8-	chr4	55152457	0+2-	DEL	342	85	2	04-.bwa.drm.sorted.bam|2	343.92
chr4	55561546	2+0-	chr4	55561547	64+38-	DEL	210	99	22	04-.bwa.drm.sorted.bam|22	2756.07
chr4	55561473	3+0-	chr4	55561547	64+38-	DEL	210	94	3	04-.bwa.drm.sorted.bam|3	2718.82
chr4	55589625	4+0-	chr4	55589636	71+71-	DEL	214	99	60	04-.bwa.drm.sorted.bam|60	2976.23
chr4	55589571	3+0-	chr4	55589636	71+71-	DEL	218	96	3	04-.bwa.drm.sorted.bam|3	5952.45
chr4	55591805	48+37-	chr4	55592190	48+37-	DEL	208	99	28	04-.bwa.drm.sorted.bam|28	NA
chr4	55592190	48+37-	chr4	55592242	0+2-	DEL	241	69	2	04-.bwa.drm.sorted.bam|2	12202.52
chr4	55593371	149+105-	chr4	55594519	149+105-	DEL	212	99	84	04-.bwa.drm.sorted.bam|84	NA
chr4	55598991	58+46-	chr4	55599570	58+46-	DEL	223	99	42	04-.bwa.drm.sorted.bam|42	NA
chr4	55599570	58+46-	chr4	55599621	0+3-	DEL	239	90	3	04-.bwa.drm.sorted.bam|3	303.46
chr4	81435107	5+0-	chr4	81435164	6+4-	DEL	186	99	4	04-.bwa.drm.sorted.bam|4	2443.64
chr4	81435288	6+4-	chr4	81435348	0+4-	DEL	187	99	3	04-.bwa.drm.sorted.bam|3	3095.27
chr4	82931630	7+0-	chr4	82931682	19+23-	DEL	238	99	22	04-.bwa.drm.sorted.bam|22	2976.23
chr4	83501420	5+1-	chr4	83501533	0+2-	DEL	167	91	2	04-.bwa.drm.sorted.bam|2	4930.53
chr4	106154782	713+518-	chr4	106158878	713+518-	DEL	212	99	453	04-.bwa.drm.sorted.bam|453	NA
chr4	106162189	11+0-	chr4	106162271	41+37-	DEL	208	99	26	04-.bwa.drm.sorted.bam|26	2076.10
chr4	106162665	41+37-	chr4	106162782	0+3-	DEL	201	99	3	04-.bwa.drm.sorted.bam|3	793.66
chr4	106163692	8+0-	chr4	106163760	59+51-	DEL	241	99	44	04-.bwa.drm.sorted.bam|44	455.19
chr4	106164336	59+51-	chr4	106164429	0+2-	DEL	370	68	2	04-.bwa.drm.sorted.bam|2	NA
chr4	106164764	47+32-	chr4	106165127	47+32-	DEL	194	99	27	04-.bwa.drm.sorted.bam|27	NA
chr4	106180582	4+0-	chr4	106180634	59+48-	DEL	203	99	39	04-.bwa.drm.sorted.bam|39	2678.60
chr4	106181190	59+48-	chr4	106181244	0+2-	DEL	359	68	2	04-.bwa.drm.sorted.bam|2	286.60
chr4	106182713	97+90-	chr4	106183222	97+90-	DEL	215	99	84	04-.bwa.drm.sorted.bam|84	NA
chr4	106190550	50+41-	chr4	106190974	50+41-	DEL	193	99	33	04-.bwa.drm.sorted.bam|33	NA
chr4	106193720	94+78-	chr4	106194195	94+78-	DEL	215	99	66	04-.bwa.drm.sorted.bam|66	NA
chr4	106195959	8+0-	chr4	106196020	160+100-	DEL	190	99	71	04-.bwa.drm.sorted.bam|71	7865.04
chr4	106197676	160+100-	chr4	106197800	0+4-	DEL	191	98	4	04-.bwa.drm.sorted.bam|4	4617.95
chr4	153245213	82+63-	chr4	153246067	82+63-	DEL	213	99	49	04-.bwa.drm.sorted.bam|49	NA
chr4	153246908	3+0-	chr4	153247031	57+14-	DEL	258	99	4	04-.bwa.drm.sorted.bam|4	2078.92
chr4	153246950	7+0-	chr4	153247031	57+14-	DEL	167	99	7	04-.bwa.drm.sorted.bam|7	3821.33
chr4	153247384	57+14-	chr4	153247448	4+34-	DEL	195	99	34	04-.bwa.drm.sorted.bam|34	4352.73
chr4	153247529	57+14-	chr4	153247698	0+3-	DEL	310	99	3	04-.bwa.drm.sorted.bam|3	11582.63
chr4	153249407	82+75-	chr4	153249922	82+75-	DEL	214	99	67	04-.bwa.drm.sorted.bam|67	NA
chr4	159336595	2+0-	chr4	159336642	0+2-	DEL	199	98	2	04-.bwa.drm.sorted.bam|2	241.82
chr5	23303621	2+0-	chr5	23303737	18+6-	DEL	194	99	4	04-.bwa.drm.sorted.bam|4	533.67
chr5	23304744	2+0-	chr5	23304817	11+3-	DEL	236	99	3	04-.bwa.drm.sorted.bam|3	780.92
chr5	23305023	11+3-	chr5	23305098	0+6-	DEL	199	99	6	04-.bwa.drm.sorted.bam|6	2888.92
chr5	93018387	61+59-	chr5	93018869	61+59-	DEL	220	99	51	04-.bwa.drm.sorted.bam|51	NA
chr5	112227269	225+171-	chr5	112228930	225+171-	DEL	218	99	149	04-.bwa.drm.sorted.bam|149	NA
chr5	170837145	5+0-	chr5	170837207	106+99-	DEL	220	99	98	04-.bwa.drm.sorted.bam|98	249.62
chr6	7517739	4+0-	chr6	7517745	11+5-	DEL	227	99	4	04-.bwa.drm.sorted.bam|4	18756.13
chr6	7518034	11+5-	chr6	7518047	0+3-	DEL	177	99	3	04-.bwa.drm.sorted.bam|3	2154.94
chr6	7517670	3+2-	chr6	7517681	3+2-	ITX	-10	99	2	04-.bwa.drm.sorted.bam|2	NA
chr6	17325513	3+0-	chr6	17325565	0+3-	DEL	213	99	3	04-.bwa.drm.sorted.bam|3	2042.57
chr6	45390421	5+0-	chr6	45390528	3+4-	DEL	208	88	2	04-.bwa.drm.sorted.bam|2	1880.31
chr6	45390566	5+0-	chr6	45390652	0+3-	DEL	174	99	3	04-.bwa.drm.sorted.bam|3	4354.82
chr6	54635306	31+22-	chr6	54635650	31+22-	DEL	185	99	15	04-.bwa.drm.sorted.bam|15	NA
chr6	54635650	31+22-	chr6	54635705	0+2-	DEL	242	70	2	04-.bwa.drm.sorted.bam|2	281.39
chr6	55804513	35+35-	chr6	55804892	35+35-	DEL	227	99	31	04-.bwa.drm.sorted.bam|31	NA
chr6	70414977	75+65-	chr6	70415334	75+65-	DEL	202	99	59	04-.bwa.drm.sorted.bam|59	NA
chr6	70415334	75+65-	chr6	70415405	0+3-	DEL	319	96	3	04-.bwa.drm.sorted.bam|3	217.98
chr6	100498038	62+31-	chr6	100498276	62+31-	DEL	206	99	28	04-.bwa.drm.sorted.bam|28	NA
chr6	100498276	62+31-	chr6	100498339	0+24-	DEL	257	99	24	04-.bwa.drm.sorted.bam|24	1473.94
chr6	138027939	6+0-	chr6	138028014	30+23-	DEL	195	99	23	04-.bwa.drm.sorted.bam|23	10523.93
chr6	138028339	30+23-	chr6	138028393	0+2-	DEL	339	75	2	04-.bwa.drm.sorted.bam|2	286.60
chr6	146726582	2+0-	chr6	146726727	0+2-	DEL	169	96	2	04-.bwa.drm.sorted.bam|2	320.20
chr7	11296966	5+0-	chr7	11297071	22+16-	DEL	209	99	13	04-.bwa.drm.sorted.bam|13	1768.73
chr7	11297333	22+16-	chr7	11297456	0+5-	DEL	235	99	5	04-.bwa.drm.sorted.bam|5	629.12
chr7	12632889	7+2-	chr7	12632965	0+2-	DEL	221	81	2	04-.bwa.drm.sorted.bam|2	2850.91
chr7	12633034	7+2-	chr7	12633064	0+3-	DEL	254	99	3	04-.bwa.drm.sorted.bam|3	1591.86
chr7	23344171	2+2-	chr7	23344223	2+2-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	47092446	2+0-	chr7	47092484	0+2-	DEL	177	93	2	04-.bwa.drm.sorted.bam|2	4905.08
chr7	50358416	88+76-	chr7	50359161	88+76-	DEL	204	99	70	04-.bwa.drm.sorted.bam|70	NA
chr7	50367203	8+0-	chr7	50367261	12+9-	DEL	165	99	5	04-.bwa.drm.sorted.bam|5	10406.53
chr7	50367374	12+9-	chr7	50367511	0+5-	DEL	205	99	5	04-.bwa.drm.sorted.bam|5	6213.14
chr7	50444132	79+55-	chr7	50444672	79+55-	DEL	197	99	40	04-.bwa.drm.sorted.bam|40	NA
chr7	50444817	79+55-	chr7	50444876	0+4-	DEL	289	99	4	04-.bwa.drm.sorted.bam|4	606.92
chr7	50449992	2+0-	chr7	50450066	16+12-	DEL	227	99	5	04-.bwa.drm.sorted.bam|5	1342.70
chr7	50454828	30+25-	chr7	50455119	30+25-	DEL	199	99	24	04-.bwa.drm.sorted.bam|24	NA
chr7	50459197	4+0-	chr7	50459262	105+92-	DEL	211	99	82	04-.bwa.drm.sorted.bam|82	9523.92
chr7	50467497	15+6-	chr7	50467661	15+6-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr7	50467806	15+6-	chr7	50467807	8+7-	DEL	210	99	4	04-.bwa.drm.sorted.bam|4	9540.23
chr7	50468051	36+11-	chr7	50468428	36+11-	ITX	-12	99	7	04-.bwa.drm.sorted.bam|7	NA
chr7	50468428	36+11-	chr7	50468542	0+10-	DEL	211	99	10	04-.bwa.drm.sorted.bam|10	6787.88
chr7	56978158	2+0-	chr7	56978261	8+5-	DEL	189	99	4	04-.bwa.drm.sorted.bam|4	1502.56
chr7	56978457	8+5-	chr7	56978531	2+2-	DEL	243	77	2	04-.bwa.drm.sorted.bam|2	5019.36
chr7	56978772	2+2-	chr7	56978856	0+2-	DEL	254	88	2	04-.bwa.drm.sorted.bam|2	608.24
chr7	57099616	5+0-	chr7	57099720	4+4-	DEL	224	99	3	04-.bwa.drm.sorted.bam|3	297.62
chr7	57099761	5+0-	chr7	57099862	0+4-	DEL	269	89	2	04-.bwa.drm.sorted.bam|2	3963.46
chr7	57099810	4+4-	chr7	57099862	0+4-	DEL	161	87	2	04-.bwa.drm.sorted.bam|2	6845.32
chr7	63005007	24+11-	chr7	63005138	24+11-	DEL	171	99	10	04-.bwa.drm.sorted.bam|10	NA
chr7	63005138	24+11-	chr7	63005197	0+9-	DEL	255	99	9	04-.bwa.drm.sorted.bam|9	262.31
chr7	63126442	20+11-	chr7	63126585	20+11-	DEL	194	99	7	04-.bwa.drm.sorted.bam|7	NA
chr7	101459289	3+0-	chr7	101459385	0+2-	DEL	175	99	2	04-.bwa.drm.sorted.bam|2	10852.72
chr7	101460796	25+8-	chr7	101461125	25+8-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr7	101461125	25+8-	chr7	101461235	0+9-	DEL	234	99	9	04-.bwa.drm.sorted.bam|9	6190.55
chr7	101559188	4+0-	chr7	101559259	38+25-	DEL	201	99	20	04-.bwa.drm.sorted.bam|20	3051.68
chr7	101671296	48+34-	chr7	101671578	48+34-	DEL	208	99	25	04-.bwa.drm.sorted.bam|25	NA
chr7	101713508	58+46-	chr7	101713944	58+46-	DEL	214	99	34	04-.bwa.drm.sorted.bam|34	NA
chr7	101740658	85+69-	chr7	101741076	85+69-	DEL	214	99	65	04-.bwa.drm.sorted.bam|65	NA
chr7	101747410	41+30-	chr7	101747855	41+30-	DEL	227	99	24	04-.bwa.drm.sorted.bam|24	NA
chr7	101747855	41+30-	chr7	101747916	0+7-	DEL	234	99	7	04-.bwa.drm.sorted.bam|7	253.71
chr7	101754719	5+0-	chr7	101755141	27+13-	ITX	-12	99	6	04-.bwa.drm.sorted.bam|6	733.48
chr7	101754996	27+13-	chr7	101755121	6+6-	DEL	224	99	4	04-.bwa.drm.sorted.bam|4	6561.98
chr7	101755211	6+6-	chr7	101755326	0+3-	DEL	180	88	2	04-.bwa.drm.sorted.bam|2	1076.62
chr7	101758172	53+39-	chr7	101758672	53+39-	DEL	219	99	37	04-.bwa.drm.sorted.bam|37	NA
chr7	101801851	48+41-	chr7	101802133	48+41-	DEL	191	99	32	04-.bwa.drm.sorted.bam|32	NA
chr7	101813470	41+27-	chr7	101813952	41+27-	DEL	201	99	23	04-.bwa.drm.sorted.bam|23	NA
chr7	101821670	37+17-	chr7	101822108	37+17-	ITX	-13	99	13	04-.bwa.drm.sorted.bam|13	NA
chr7	101822108	37+17-	chr7	101822221	0+6-	DEL	202	99	6	04-.bwa.drm.sorted.bam|6	8902.34
chr7	101833096	22+8-	chr7	101833177	22+8-	DEL	167	99	3	04-.bwa.drm.sorted.bam|3	NA
chr7	101833177	22+8-	chr7	101833253	2+3-	DEL	198	79	2	04-.bwa.drm.sorted.bam|2	7941.82
chr7	101836959	2+0-	chr7	101837100	31+6-	DEL	166	99	5	04-.bwa.drm.sorted.bam|5	8341.87
chr7	101837296	31+6-	chr7	101837360	0+25-	DEL	241	99	24	04-.bwa.drm.sorted.bam|24	6770.91
chr7	101838712	12+7-	chr7	101838900	12+7-	ITX	-12	99	5	04-.bwa.drm.sorted.bam|5	NA
chr7	101838900	12+7-	chr7	101839020	0+3-	DEL	176	99	3	04-.bwa.drm.sorted.bam|3	10059.64
chr7	101839722	89+57-	chr7	101840527	89+57-	DEL	198	99	44	04-.bwa.drm.sorted.bam|44	NA
chr7	101840527	89+57-	chr7	101840596	3+4-	DEL	177	86	3	04-.bwa.drm.sorted.bam|3	10093.29
chr7	101841947	38+27-	chr7	101842416	38+27-	DEL	184	99	20	04-.bwa.drm.sorted.bam|20	NA
chr7	101843033	4+0-	chr7	101843090	50+40-	DEL	201	99	34	04-.bwa.drm.sorted.bam|34	271.52
chr7	101843646	50+40-	chr7	101843714	0+2-	DEL	260	68	2	04-.bwa.drm.sorted.bam|2	910.37
chr7	101844444	2+0-	chr7	101844503	10+4-	DEL	176	99	3	04-.bwa.drm.sorted.bam|3	4196.98
chr7	101844688	10+4-	chr7	101844739	7+5-	DEL	162	99	4	04-.bwa.drm.sorted.bam|4	19117.87
chr7	101844847	7+5-	chr7	101844911	49+22-	DEL	166	99	12	04-.bwa.drm.sorted.bam|12	15476.37
chr7	101845653	49+22-	chr7	101845773	0+2-	DEL	262	65	2	04-.bwa.drm.sorted.bam|2	1547.64
chr7	101847542	10+3-	chr7	101847731	10+3-	ITX	-10	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	101848194	5+0-	chr7	101848272	23+18-	DEL	208	99	11	04-.bwa.drm.sorted.bam|11	2845.43
chr7	101848270	2+0-	chr7	101848272	23+18-	DEL	168	74	2	04-.bwa.drm.sorted.bam|2	4105.98
chr7	101870413	12+0-	chr7	101870469	32+33-	DEL	213	99	26	04-.bwa.drm.sorted.bam|26	1934.55
chr7	101877279	3+0-	chr7	101877283	33+23-	DEL	188	99	14	04-.bwa.drm.sorted.bam|14	9036.54
chr7	101877668	33+23-	chr7	101877798	0+4-	DEL	222	99	4	04-.bwa.drm.sorted.bam|4	5119.11
chr7	101882662	34+17-	chr7	101882980	34+17-	DEL	190	99	9	04-.bwa.drm.sorted.bam|9	NA
chr7	101882980	34+17-	chr7	101883031	0+2-	DEL	187	71	2	04-.bwa.drm.sorted.bam|2	19117.87
chr7	101882980	34+17-	chr7	101883117	0+2-	DEL	195	71	2	04-.bwa.drm.sorted.bam|2	10957.72
chr7	101883125	34+17-	chr7	101883176	0+2-	DEL	184	71	2	04-.bwa.drm.sorted.bam|2	7817.15
chr7	101916648	15+6-	chr7	101916812	15+6-	DEL	179	99	3	04-.bwa.drm.sorted.bam|3	NA
chr7	101916812	15+6-	chr7	101916946	0+2-	DEL	159	75	2	04-.bwa.drm.sorted.bam|2	4157.83
chr7	101917384	7+2-	chr7	101917457	7+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	101917457	7+2-	chr7	101917530	13+5-	DEL	181	99	3	04-.bwa.drm.sorted.bam|3	9752.23
chr7	101918490	18+3-	chr7	101918662	18+3-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	101921219	4+3-	chr7	101921267	4+3-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	101923210	14+8-	chr7	101923539	14+8-	DEL	194	99	7	04-.bwa.drm.sorted.bam|7	NA
chr7	101923947	7+4-	chr7	101924040	7+4-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	NA
chr7	101924117	13+7-	chr7	101924375	13+7-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	NA
chr7	101925051	3+2-	chr7	101925108	3+2-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chr7	112161472	12+0-	chr7	112161560	10+10-	DEL	189	99	10	04-.bwa.drm.sorted.bam|10	175.87
chr7	112161617	12+0-	chr7	112161781	0+6-	DEL	337	99	3	04-.bwa.drm.sorted.bam|3	4357.42
chr7	112161726	10+10-	chr7	112161781	0+6-	DEL	184	99	3	04-.bwa.drm.sorted.bam|3	844.17
chr7	112161871	10+10-	chr7	112161909	0+2-	DEL	229	84	2	04-.bwa.drm.sorted.bam|2	845.70
chr7	117962499	2+1-	chr7	117962541	0+2-	DEL	221	91	2	04-.bwa.drm.sorted.bam|2	165.52
chr7	140452870	24+0-	chr7	140452950	33+50-	DEL	232	99	43	04-.bwa.drm.sorted.bam|43	4062.55
chr7	148504574	41+41-	chr7	148504957	41+41-	DEL	213	99	34	04-.bwa.drm.sorted.bam|34	NA
chr7	148505981	86+65-	chr7	148506718	86+65-	DEL	217	99	60	04-.bwa.drm.sorted.bam|60	NA
chr7	148507385	36+25-	chr7	148507682	36+25-	DEL	183	99	21	04-.bwa.drm.sorted.bam|21	NA
chr7	148508641	22+18-	chr7	148508987	22+18-	DEL	213	99	15	04-.bwa.drm.sorted.bam|15	NA
chr7	148510818	6+0-	chr7	148510882	27+14-	DEL	184	99	10	04-.bwa.drm.sorted.bam|10	12090.92
chr7	148511275	27+14-	chr7	148511348	0+2-	DEL	190	73	2	04-.bwa.drm.sorted.bam|2	2332.06
chr7	148511635	3+0-	chr7	148511693	94+66-	DEL	211	99	53	04-.bwa.drm.sorted.bam|53	266.83
chr7	148512791	94+66-	chr7	148512849	0+2-	DEL	262	60	2	04-.bwa.drm.sorted.bam|2	1601.00
chr7	148512936	94+66-	chr7	148513003	0+2-	DEL	347	60	2	04-.bwa.drm.sorted.bam|2	803.02
chr7	148513507	10+0-	chr7	148513559	234+208-	DEL	213	99	181	04-.bwa.drm.sorted.bam|181	595.25
chr7	148516406	2+0-	chr7	148516526	65+51-	DEL	219	99	49	04-.bwa.drm.sorted.bam|49	773.82
chr7	148523337	166+148-	chr7	148524573	166+148-	DEL	217	99	137	04-.bwa.drm.sorted.bam|137	NA
chr7	148525517	5+0-	chr7	148525568	72+62-	DEL	219	99	49	04-.bwa.drm.sorted.bam|49	303.46
chr7	148526479	6+0-	chr7	148526531	84+76-	DEL	214	99	70	04-.bwa.drm.sorted.bam|70	297.62
chr7	148527177	84+76-	chr7	148527247	0+2-	DEL	253	66	2	04-.bwa.drm.sorted.bam|2	221.09
chr7	148529595	42+32-	chr7	148530070	42+32-	DEL	209	99	27	04-.bwa.drm.sorted.bam|27	NA
chr7	148543276	7+0-	chr7	148543376	74+61-	DEL	200	99	52	04-.bwa.drm.sorted.bam|52	2785.75
chr7	148543846	74+61-	chr7	148543914	90+51-	DEL	207	99	46	04-.bwa.drm.sorted.bam|46	455.19
chr7	148544429	90+51-	chr7	148544480	0+21-	DEL	207	99	21	04-.bwa.drm.sorted.bam|21	8496.83
chr7	149031591	8+0-	chr7	149031649	58+59-	DEL	239	99	56	04-.bwa.drm.sorted.bam|56	266.83
chr7	153442559	3+0-	chr7	153442703	6+8-	DEL	207	99	6	04-.bwa.drm.sorted.bam|6	429.90
chr8	48649832	4+0-	chr8	48649958	3+2-	DEL	165	87	2	04-.bwa.drm.sorted.bam|2	4053.34
chr8	48649977	4+0-	chr8	48650083	0+2-	DEL	199	87	2	04-.bwa.drm.sorted.bam|2	7645.70
chr8	59338378	2+0-	chr8	59338446	4+3-	DEL	185	86	2	04-.bwa.drm.sorted.bam|2	1820.75
chr8	59338727	4+3-	chr8	59338752	0+2-	DEL	195	86	2	04-.bwa.drm.sorted.bam|2	3732.54
chr8	59338903	2+0-	chr8	59338954	5+3-	DEL	166	84	2	04-.bwa.drm.sorted.bam|2	303.46
chr8	62115484	71+56-	chr8	62115893	71+56-	DEL	218	99	54	04-.bwa.drm.sorted.bam|54	NA
chr8	62115893	71+56-	chr8	62116024	0+3-	DEL	338	95	3	04-.bwa.drm.sorted.bam|3	1063.26
chr8	68098113	63+56-	chr8	68098452	63+56-	DEL	216	99	50	04-.bwa.drm.sorted.bam|50	NA
chr8	117859554	10+0-	chr8	117859624	58+52-	DEL	194	99	45	04-.bwa.drm.sorted.bam|45	2653.09
chr8	117860891	138+124-	chr8	117861481	138+124-	DEL	213	99	117	04-.bwa.drm.sorted.bam|117	NA
chr8	117862616	97+88-	chr8	117863297	97+88-	DEL	222	99	80	04-.bwa.drm.sorted.bam|80	NA
chr8	117864060	8+0-	chr8	117864115	25+13-	DEL	180	99	9	04-.bwa.drm.sorted.bam|9	16601.93
chr8	117864320	25+13-	chr8	117864378	2+7-	DEL	203	99	7	04-.bwa.drm.sorted.bam|7	2668.34
chr8	117864465	25+13-	chr8	117864504	59+50-	DEL	206	99	43	04-.bwa.drm.sorted.bam|43	2018.66
chr8	117864438	2+7-	chr8	117864504	59+50-	DEL	301	65	2	04-.bwa.drm.sorted.bam|2	234.49
chr8	117866174	112+91-	chr8	117866888	112+91-	DEL	216	99	84	04-.bwa.drm.sorted.bam|84	NA
chr8	117868267	2+0-	chr8	117868314	18+4-	DEL	226	88	2	04-.bwa.drm.sorted.bam|2	2901.82
chr8	117868406	18+4-	chr8	117868509	8+6-	DEL	196	99	6	04-.bwa.drm.sorted.bam|6	4507.68
chr8	117868702	8+6-	chr8	117868764	180+166-	DEL	222	99	156	04-.bwa.drm.sorted.bam|156	6739.71
chr8	117870232	11+0-	chr8	117870288	93+82-	DEL	211	99	72	04-.bwa.drm.sorted.bam|72	2763.64
chr8	117873872	4+0-	chr8	117873936	54+51-	DEL	207	99	39	04-.bwa.drm.sorted.bam|39	1110.74
chr8	117873872	10+0-	chr8	117873936	54+51-	DEL	216	99	10	04-.bwa.drm.sorted.bam|10	725.45
chr8	117874359	54+51-	chr8	117874412	0+2-	DEL	253	72	2	04-.bwa.drm.sorted.bam|2	292.01
chr8	117874359	54+51-	chr8	117874484	0+2-	DEL	246	71	2	04-.bwa.drm.sorted.bam|2	371.43
chr8	117875196	63+49-	chr8	117875730	63+49-	DEL	222	99	44	04-.bwa.drm.sorted.bam|44	NA
chr8	117878463	3+0-	chr8	117878522	68+62-	DEL	239	99	61	04-.bwa.drm.sorted.bam|61	262.31
chr8	117879234	68+62-	chr8	117879288	0+3-	DEL	425	89	3	04-.bwa.drm.sorted.bam|3	NA
chr8	129255236	3+0-	chr8	129255329	1+2-	DEL	159	89	2	04-.bwa.drm.sorted.bam|2	1164.89
chr9	5069617	2+0-	chr9	5069731	103+103-	DEL	233	99	86	04-.bwa.drm.sorted.bam|86	1374.35
chr9	5069677	13+0-	chr9	5069731	103+103-	DEL	235	99	13	04-.bwa.drm.sorted.bam|13	2865.99
chr9	5073415	4+0-	chr9	5073477	64+55-	DEL	212	99	53	04-.bwa.drm.sorted.bam|53	1248.09
chr9	21968242	16+5-	chr9	21968382	56+58-	DEL	203	99	53	04-.bwa.drm.sorted.bam|53	11938.92
chr9	21968331	2+1-	chr9	21968382	56+58-	DEL	171	66	2	04-.bwa.drm.sorted.bam|2	14869.45
chr9	21970651	2+0-	chr9	21970776	6+3-	DEL	167	92	2	04-.bwa.drm.sorted.bam|2	1733.35
chr9	21970847	6+3-	chr9	21970929	2+4-	DEL	178	99	3	04-.bwa.drm.sorted.bam|3	3963.46
chr9	21970992	6+3-	chr9	21971064	1+2-	DEL	185	89	2	04-.bwa.drm.sorted.bam|2	5135.02
chr9	21974146	24+13-	chr9	21974556	24+13-	ITX	-12	99	7	04-.bwa.drm.sorted.bam|7	NA
chr9	21974556	24+13-	chr9	21974621	2+2-	DEL	235	72	2	04-.bwa.drm.sorted.bam|2	4047.67
chr9	21974810	2+2-	chr9	21974960	0+4-	DEL	237	97	2	04-.bwa.drm.sorted.bam|2	7659.49
chr9	21994100	5+0-	chr9	21994216	5+5-	DEL	189	99	4	04-.bwa.drm.sorted.bam|4	5336.68
chr9	33675610	4+0-	chr9	33675698	20+8-	DEL	213	99	4	04-.bwa.drm.sorted.bam|4	1758.68
chr9	33675816	20+8-	chr9	33675879	78+61-	DEL	197	99	51	04-.bwa.drm.sorted.bam|51	15476.37
chr9	33676457	78+61-	chr9	33676509	0+9-	DEL	236	99	9	04-.bwa.drm.sorted.bam|9	595.25
chr9	133738035	11+1-	chr9	133738093	38+35-	DEL	206	99	27	04-.bwa.drm.sorted.bam|27	14409.04
chr9	133747248	8+0-	chr9	133747325	30+23-	DEL	205	99	17	04-.bwa.drm.sorted.bam|17	4220.83
chr9	133747649	30+23-	chr9	133747780	0+3-	DEL	178	99	3	04-.bwa.drm.sorted.bam|3	3426.07
chr9	133748084	16+7-	chr9	133748306	16+7-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr9	133748306	16+7-	chr9	133748359	3+2-	DEL	197	80	2	04-.bwa.drm.sorted.bam|2	16936.41
chr9	133748306	16+7-	chr9	133748434	1+3-	DEL	247	99	3	04-.bwa.drm.sorted.bam|3	12937.28
chr9	139390286	2+0-	chr9	139390367	6+5-	DEL	173	85	2	04-.bwa.drm.sorted.bam|2	2101.73
chr9	139390657	2+1-	chr9	139390743	38+22-	DEL	190	99	12	04-.bwa.drm.sorted.bam|12	6118.57
chr9	139391250	38+22-	chr9	139391321	42+23-	DEL	191	99	12	04-.bwa.drm.sorted.bam|12	15476.37
chr9	139391894	42+23-	chr9	139391995	0+2-	DEL	169	68	2	04-.bwa.drm.sorted.bam|2	5976.02
chr9	139396840	5+2-	chr9	139396902	19+10-	DEL	172	99	6	04-.bwa.drm.sorted.bam|6	7738.19
chr9	139397191	19+10-	chr9	139397259	1+6-	DEL	239	99	6	04-.bwa.drm.sorted.bam|6	1820.75
chr9	139397579	20+8-	chr9	139397834	20+8-	ITX	-13	99	5	04-.bwa.drm.sorted.bam|5	NA
chr9	139397834	20+8-	chr9	139397903	0+2-	DEL	178	77	2	04-.bwa.drm.sorted.bam|2	7177.45
chr9	139399148	2+2-	chr9	139399199	6+6-	DEL	203	84	2	04-.bwa.drm.sorted.bam|2	7106.50
chr9	139399123	5+2-	chr9	139399199	6+6-	DEL	180	83	2	04-.bwa.drm.sorted.bam|2	8960.00
chr10	21402492	16+17-	chr10	21402560	16+17-	DEL	163	99	6	04-.bwa.drm.sorted.bam|6	NA
chr10	74677016	3+0-	chr10	74677085	72+65-	DEL	217	99	59	04-.bwa.drm.sorted.bam|59	224.30
chr10	89692571	100+86-	chr10	89693110	100+86-	DEL	213	99	83	04-.bwa.drm.sorted.bam|83	NA
chr10	89693110	100+86-	chr10	89693163	0+6-	DEL	288	99	6	04-.bwa.drm.sorted.bam|6	876.02
chr10	89717356	111+85-	chr10	89717984	111+85-	DEL	215	99	75	04-.bwa.drm.sorted.bam|75	NA
chr10	89717984	111+85-	chr10	89718095	0+13-	DEL	229	99	13	04-.bwa.drm.sorted.bam|13	139.43
chr10	97948993	31+13-	chr10	97949126	31+13-	DEL	193	99	5	04-.bwa.drm.sorted.bam|5	NA
chr10	97949126	31+13-	chr10	97949178	0+15-	DEL	219	99	15	04-.bwa.drm.sorted.bam|15	2380.98
chr10	112341933	4+0-	chr10	112342020	101+95-	DEL	212	99	91	04-.bwa.drm.sorted.bam|91	177.89
chr10	112343818	57+45-	chr10	112344225	57+45-	DEL	205	99	43	04-.bwa.drm.sorted.bam|43	NA
chr10	112344225	57+45-	chr10	112344284	0+4-	DEL	177	99	4	04-.bwa.drm.sorted.bam|4	524.62
chr10	112355966	26+0-	chr10	112356033	53+66-	DEL	231	99	66	04-.bwa.drm.sorted.bam|66	1154.95
chr10	112356527	53+66-	chr10	112356588	0+4-	DEL	346	99	4	04-.bwa.drm.sorted.bam|4	NA
chr10	112360587	22+0-	chr10	112360642	52+72-	DEL	220	99	69	04-.bwa.drm.sorted.bam|69	2251.11
chr10	112361586	83+72-	chr10	112362010	83+72-	DEL	212	99	66	04-.bwa.drm.sorted.bam|66	NA
chr10	112362752	82+76-	chr10	112363255	82+76-	DEL	226	99	71	04-.bwa.drm.sorted.bam|71	NA
chr10	112363255	82+76-	chr10	112363340	0+2-	DEL	212	67	2	04-.bwa.drm.sorted.bam|2	182.07
chr11	533832	9+3-	chr11	533973	9+3-	ITX	-13	99	3	04-.bwa.drm.sorted.bam|3	NA
chr11	534026	4+5-	chr11	534157	4+5-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr11	32413290	8+0-	chr11	32413377	31+25-	DEL	198	99	14	04-.bwa.drm.sorted.bam|14	6759.79
chr11	32413728	31+25-	chr11	32413791	0+3-	DEL	167	99	3	04-.bwa.drm.sorted.bam|3	4667.48
chr11	32417785	4+0-	chr11	32417790	13+8-	DEL	187	99	4	04-.bwa.drm.sorted.bam|4	15063.67
chr11	32417713	7+3-	chr11	32418182	13+8-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	1649.93
chr11	32418037	13+8-	chr11	32418148	0+3-	DEL	201	99	3	04-.bwa.drm.sorted.bam|3	557.71
chr11	62099077	57+47-	chr11	62099486	57+47-	DEL	209	99	44	04-.bwa.drm.sorted.bam|44	NA
chr11	62099486	57+47-	chr11	62099539	0+3-	DEL	326	94	3	04-.bwa.drm.sorted.bam|3	292.01
chr11	71991150	6+0-	chr11	71991151	6+11-	DEL	188	99	6	04-.bwa.drm.sorted.bam|6	1484.04
chr11	74789878	5+0-	chr11	74789950	77+55-	DEL	205	99	46	04-.bwa.drm.sorted.bam|46	214.95
chr11	74790403	77+55-	chr11	74790465	0+21-	DEL	249	99	21	04-.bwa.drm.sorted.bam|21	499.24
chr11	94770797	5+2-	chr11	94770936	0+2-	DEL	170	87	2	04-.bwa.drm.sorted.bam|2	2672.18
chr11	104552816	53+42-	chr11	104553288	53+42-	DEL	226	99	37	04-.bwa.drm.sorted.bam|37	NA
chr11	104553288	53+42-	chr11	104553408	0+2-	DEL	345	67	2	04-.bwa.drm.sorted.bam|2	128.97
chr11	109345726	4+0-	chr11	109345732	1+3-	DEL	204	99	3	04-.bwa.drm.sorted.bam|3	922.43
chr11	118326907	0+20-	chr11	118354267	893+713-	DEL	211	99	607	04-.bwa.drm.sorted.bam|607	17635.36
chr11	118354213	19+0-	chr11	118354267	893+713-	DEL	191	99	19	04-.bwa.drm.sorted.bam|19	7164.99
chr11	118358567	893+713-	chr11	118358621	95+83-	DEL	205	99	68	04-.bwa.drm.sorted.bam|68	3725.79
chr11	118359586	95+83-	chr11	118359731	2+3-	DEL	186	85	3	04-.bwa.drm.sorted.bam|3	2027.94
chr11	118359812	2+3-	chr11	118359872	190+153-	DEL	206	99	132	04-.bwa.drm.sorted.bam|132	1805.58
chr11	118361079	190+153-	chr11	118361144	0+2-	DEL	239	59	2	04-.bwa.drm.sorted.bam|2	476.20
chr11	118339368	51+34-	chr11	118339670	51+34-	DEL	211	99	30	04-.bwa.drm.sorted.bam|30	NA
chr11	118339670	51+34-	chr11	118339731	1965+1609-	DEL	212	99	1455	04-.bwa.drm.sorted.bam|1455	4313.09
chr11	118348151	1965+1609-	chr11	118348214	697+574-	DEL	211	99	513	04-.bwa.drm.sorted.bam|513	736.97
chr11	118351122	697+574-	chr11	118351257	0+5-	DEL	281	99	5	04-.bwa.drm.sorted.bam|5	1031.76
chr11	118352281	230+162-	chr11	118353621	230+162-	DEL	216	99	147	04-.bwa.drm.sorted.bam|147	NA
chr11	118353621	230+162-	chr11	118353672	13+14-	DEL	181	99	12	04-.bwa.drm.sorted.bam|12	7586.46
chr11	118353766	230+162-	chr11	118353933	1+10-	DEL	278	55	2	04-.bwa.drm.sorted.bam|2	10168.77
chr11	118353873	13+14-	chr11	118353933	1+10-	DEL	211	99	8	04-.bwa.drm.sorted.bam|8	5674.67
chr11	118373766	88+74-	chr11	118374421	88+74-	DEL	218	99	67	04-.bwa.drm.sorted.bam|67	NA
chr11	119148673	24+15-	chr11	119148851	24+15-	DEL	198	99	13	04-.bwa.drm.sorted.bam|13	NA
chr11	119148851	24+15-	chr11	119148906	93+77-	DEL	225	99	60	04-.bwa.drm.sorted.bam|60	11536.93
chr11	119328842	3+1-	chr11	119328976	0+3-	DEL	205	99	3	04-.bwa.drm.sorted.bam|3	230.99
chr12	9848549	85+71-	chr12	9848984	85+71-	DEL	222	99	67	04-.bwa.drm.sorted.bam|67	NA
chr12	11803081	9+3-	chr12	11803178	9+3-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr12	11905526	12+1-	chr12	11905549	3+4-	DEL	210	99	3	04-.bwa.drm.sorted.bam|3	8475.16
chr12	11991971	60+47-	chr12	11992477	60+47-	DEL	216	99	40	04-.bwa.drm.sorted.bam|40	NA
chr12	11992477	60+47-	chr12	11992547	0+2-	DEL	354	66	2	04-.bwa.drm.sorted.bam|2	442.18
chr12	12006191	60+38-	chr12	12006690	60+38-	DEL	223	99	33	04-.bwa.drm.sorted.bam|33	NA
chr12	12022298	4+0-	chr12	12022366	32+19-	DEL	207	99	9	04-.bwa.drm.sorted.bam|9	7483.88
chr12	12022898	32+19-	chr12	12023022	0+6-	DEL	214	99	6	04-.bwa.drm.sorted.bam|6	4617.95
chr12	12023043	32+19-	chr12	12023162	0+2-	DEL	293	69	2	04-.bwa.drm.sorted.bam|2	2579.40
chr12	12037100	4+0-	chr12	12037164	60+53-	DEL	201	99	48	04-.bwa.drm.sorted.bam|48	5561.82
chr12	12038696	49+36-	chr12	12039214	49+36-	DEL	204	99	34	04-.bwa.drm.sorted.bam|34	NA
chr12	12039214	49+36-	chr12	12039275	0+2-	DEL	263	67	2	04-.bwa.drm.sorted.bam|2	253.71
chr12	12043690	45+24-	chr12	12044120	45+24-	DEL	202	99	20	04-.bwa.drm.sorted.bam|20	NA
chr12	12044120	45+24-	chr12	12044227	0+3-	DEL	181	94	3	04-.bwa.drm.sorted.bam|3	1735.67
chr12	25379829	3+0-	chr12	25379893	68+62-	DEL	211	99	52	04-.bwa.drm.sorted.bam|52	241.82
chr12	25398068	74+60-	chr12	25398606	74+60-	DEL	206	99	49	04-.bwa.drm.sorted.bam|49	NA
chr12	49748038	3+2-	chr12	49748074	3+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr12	112887855	4+0-	chr12	112887917	60+37-	DEL	194	99	24	04-.bwa.drm.sorted.bam|24	1996.95
chr12	112888469	60+37-	chr12	112888553	0+4-	DEL	178	99	4	04-.bwa.drm.sorted.bam|4	1658.18
chr12	112888614	60+37-	chr12	112888689	0+2-	DEL	250	69	2	04-.bwa.drm.sorted.bam|2	984.86
chr12	112926580	8+0-	chr12	112926677	26+22-	DEL	184	99	13	04-.bwa.drm.sorted.bam|13	4148.31
chr12	112927037	26+22-	chr12	112927159	0+3-	DEL	223	99	3	04-.bwa.drm.sorted.bam|3	1141.70
chr13	19455806	4+0-	chr13	19455861	20+15-	DEL	204	99	12	04-.bwa.drm.sorted.bam|12	844.17
chr13	19459226	7+0-	chr13	19459294	12+12-	DEL	222	99	10	04-.bwa.drm.sorted.bam|10	910.37
chr13	19459535	12+12-	chr13	19459651	0+3-	DEL	206	99	3	04-.bwa.drm.sorted.bam|3	3602.26
chr13	19626711	15+7-	chr13	19626860	15+7-	DEL	208	99	5	04-.bwa.drm.sorted.bam|5	NA
chr13	19626860	15+7-	chr13	19626941	0+3-	DEL	175	99	3	04-.bwa.drm.sorted.bam|3	2674.93
chr13	19943480	39+33-	chr13	19943742	39+33-	DEL	190	99	33	04-.bwa.drm.sorted.bam|33	NA
chr13	20508568	22+0-	chr13	20508633	16+36-	DEL	201	99	34	04-.bwa.drm.sorted.bam|34	7381.04
chr13	20867018	3+0-	chr13	20867040	7+5-	DEL	214	99	3	04-.bwa.drm.sorted.bam|3	4262.95
chr13	20867127	7+5-	chr13	20867262	0+3-	DEL	170	99	3	04-.bwa.drm.sorted.bam|3	9285.82
chr13	20877432	2+0-	chr13	20877989	13+11-	ITX	-13	99	6	04-.bwa.drm.sorted.bam|6	944.70
chr13	20877628	2+0-	chr13	20877688	13+11-	DEL	211	82	2	04-.bwa.drm.sorted.bam|2	6190.55
chr13	21667148	17+0-	chr13	21667229	8+22-	DEL	214	99	17	04-.bwa.drm.sorted.bam|17	1719.60
chr13	21686893	6+2-	chr13	21686929	6+2-	ITX	-10	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	22520627	6+0-	chr13	22520741	11+10-	DEL	188	99	6	04-.bwa.drm.sorted.bam|6	1221.82
chr13	22605450	5+0-	chr13	22605472	6+7-	DEL	192	99	4	04-.bwa.drm.sorted.bam|4	2965.53
chr13	22606105	6+0-	chr13	22606189	15+8-	DEL	183	99	6	04-.bwa.drm.sorted.bam|6	1289.70
chr13	22606297	15+8-	chr13	22606377	3+11-	DEL	199	99	10	04-.bwa.drm.sorted.bam|10	8898.91
chr13	22731084	13+6-	chr13	22731270	13+6-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	22731415	13+6-	chr13	22731472	0+4-	DEL	260	99	4	04-.bwa.drm.sorted.bam|4	2298.47
chr13	23427397	3+0-	chr13	23427505	46+42-	DEL	229	99	40	04-.bwa.drm.sorted.bam|40	143.30
chr13	23515436	22+21-	chr13	23515709	22+21-	DEL	213	99	20	04-.bwa.drm.sorted.bam|20	NA
chr13	23553404	12+3-	chr13	23553510	12+3-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	23553510	12+3-	chr13	23553566	0+2-	DEL	155	89	2	04-.bwa.drm.sorted.bam|2	4421.82
chr13	23553510	12+3-	chr13	23553630	0+2-	DEL	175	87	2	04-.bwa.drm.sorted.bam|2	3998.06
chr13	23965912	3+0-	chr13	23966001	11+4-	DEL	182	99	3	04-.bwa.drm.sorted.bam|3	4173.40
chr13	24012773	4+0-	chr13	24012854	6+3-	DEL	174	88	2	04-.bwa.drm.sorted.bam|2	4394.52
chr13	24012918	4+0-	chr13	24013030	0+3-	DEL	238	95	2	04-.bwa.drm.sorted.bam|2	5058.42
chr13	24275367	9+5-	chr13	24275549	9+5-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	24275549	9+5-	chr13	24275631	0+6-	DEL	191	99	6	04-.bwa.drm.sorted.bam|6	2076.10
chr13	24541213	15+0-	chr13	24541296	13+12-	DEL	193	99	9	04-.bwa.drm.sorted.bam|9	3915.71
chr13	24541358	15+0-	chr13	24541477	0+10-	DEL	295	99	5	04-.bwa.drm.sorted.bam|5	13014.22
chr13	24541421	13+12-	chr13	24541477	0+10-	DEL	183	99	5	04-.bwa.drm.sorted.bam|5	9396.37
chr13	24817862	18+13-	chr13	24818114	18+13-	DEL	199	99	10	04-.bwa.drm.sorted.bam|10	NA
chr13	24937160	20+0-	chr13	24937227	6+21-	DEL	199	99	18	04-.bwa.drm.sorted.bam|18	14321.42
chr13	24937305	20+0-	chr13	24937442	0+5-	DEL	205	83	2	04-.bwa.drm.sorted.bam|2	13281.14
chr13	24937378	6+21-	chr13	24937442	0+5-	DEL	180	99	3	04-.bwa.drm.sorted.bam|3	1934.55
chr13	25035095	12+0-	chr13	25035149	14+15-	DEL	198	99	11	04-.bwa.drm.sorted.bam|11	10604.18
chr13	25035277	14+15-	chr13	25035342	0+5-	DEL	181	99	4	04-.bwa.drm.sorted.bam|4	4285.76
chr13	25049453	2+0-	chr13	25049516	87+83-	DEL	208	99	82	04-.bwa.drm.sorted.bam|82	245.66
chr13	25067236	4+0-	chr13	25067262	9+6-	DEL	223	99	5	04-.bwa.drm.sorted.bam|5	3348.69
chr13	25067590	9+6-	chr13	25067601	0+3-	DEL	235	99	3	04-.bwa.drm.sorted.bam|3	1587.32
chr13	25234902	15+2-	chr13	25235012	0+6-	DEL	191	99	6	04-.bwa.drm.sorted.bam|6	4783.61
chr13	25466870	35+33-	chr13	25467229	35+33-	DEL	200	99	31	04-.bwa.drm.sorted.bam|31	NA
chr13	25474611	9+0-	chr13	25474694	15+13-	DEL	188	99	9	04-.bwa.drm.sorted.bam|9	4475.10
chr13	25474863	15+13-	chr13	25474990	0+3-	DEL	164	99	3	04-.bwa.drm.sorted.bam|3	3046.53
chr13	25713354	3+0-	chr13	25713408	5+6-	DEL	228	99	3	04-.bwa.drm.sorted.bam|3	1088.79
chr13	26264127	33+0-	chr13	26264184	2+31-	DEL	257	99	31	04-.bwa.drm.sorted.bam|31	6787.88
chr13	26264272	33+0-	chr13	26264454	0+4-	DEL	443	74	2	04-.bwa.drm.sorted.bam|2	11595.45
chr13	26264380	2+31-	chr13	26264454	0+4-	DEL	212	79	2	04-.bwa.drm.sorted.bam|2	836.56
chr13	26307681	15+0-	chr13	26307747	16+20-	DEL	210	99	16	04-.bwa.drm.sorted.bam|16	1641.43
chr13	26307969	16+20-	chr13	26308063	0+4-	DEL	214	99	4	04-.bwa.drm.sorted.bam|4	1811.06
chr13	27402991	3+0-	chr13	27403016	8+10-	DEL	210	99	3	04-.bwa.drm.sorted.bam|3	1001.41
chr13	27402935	4+0-	chr13	27403016	8+10-	DEL	231	99	3	04-.bwa.drm.sorted.bam|3	955.33
chr13	27693008	15+4-	chr13	27693103	15+4-	DEL	194	80	2	04-.bwa.drm.sorted.bam|2	NA
chr13	27693103	15+4-	chr13	27693165	0+4-	DEL	211	99	4	04-.bwa.drm.sorted.bam|4	2246.57
chr13	28011680	2+0-	chr13	28011737	33+15-	DEL	192	99	7	04-.bwa.drm.sorted.bam|7	271.52
chr13	28011975	33+15-	chr13	28012108	0+13-	DEL	238	99	13	04-.bwa.drm.sorted.bam|13	3607.27
chr13	28270179	7+0-	chr13	28270241	51+50-	DEL	228	99	47	04-.bwa.drm.sorted.bam|47	499.24
chr13	28270736	51+50-	chr13	28270814	0+4-	DEL	433	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	28299786	10+2-	chr13	28299879	0+8-	DEL	177	99	8	04-.bwa.drm.sorted.bam|8	1996.95
chr13	28577422	148+110-	chr13	28578268	148+110-	DEL	212	99	96	04-.bwa.drm.sorted.bam|96	NA
chr13	28578268	148+110-	chr13	28578336	0+5-	DEL	231	99	5	04-.bwa.drm.sorted.bam|5	5007.06
chr13	28588413	64+55-	chr13	28588929	64+55-	DEL	201	99	52	04-.bwa.drm.sorted.bam|52	NA
chr13	28588996	3+0-	chr13	28589065	40+36-	DEL	194	99	31	04-.bwa.drm.sorted.bam|31	224.30
chr13	28589535	40+36-	chr13	28589609	2+2-	DEL	165	69	2	04-.bwa.drm.sorted.bam|2	1254.84
chr13	28592367	32+25-	chr13	28592726	32+25-	DEL	208	99	22	04-.bwa.drm.sorted.bam|22	NA
chr13	28597268	127+116-	chr13	28597750	127+116-	DEL	208	99	107	04-.bwa.drm.sorted.bam|107	NA
chr13	28598723	72+68-	chr13	28599329	72+68-	DEL	232	99	66	04-.bwa.drm.sorted.bam|66	NA
chr13	28599791	7+4-	chr13	28599888	7+4-	ITX	-14	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	28600033	7+4-	chr13	28600083	0+2-	DEL	187	88	2	04-.bwa.drm.sorted.bam|2	634.93
chr13	28601119	56+44-	chr13	28601478	56+44-	DEL	190	99	37	04-.bwa.drm.sorted.bam|37	NA
chr13	28601478	56+44-	chr13	28601570	0+3-	DEL	281	96	3	04-.bwa.drm.sorted.bam|3	504.66
chr13	28602292	43+42-	chr13	28602658	43+42-	DEL	209	99	35	04-.bwa.drm.sorted.bam|35	NA
chr13	28607658	32+2-	chr13	28607768	32+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	28607768	32+2-	chr13	28607832	111+107-	DEL	211	99	92	04-.bwa.drm.sorted.bam|92	24907.29
chr13	28609390	3+0-	chr13	28609516	17+9-	DEL	311	99	4	04-.bwa.drm.sorted.bam|4	913.73
chr13	28609722	17+9-	chr13	28609777	29+29-	DEL	190	99	28	04-.bwa.drm.sorted.bam|28	5627.77
chr13	28611142	49+40-	chr13	28611477	49+40-	DEL	195	99	38	04-.bwa.drm.sorted.bam|38	NA
chr13	28613069	7+0-	chr13	28613124	16+9-	DEL	172	99	6	04-.bwa.drm.sorted.bam|6	8441.66
chr13	28613265	16+9-	chr13	28613384	0+8-	DEL	178	99	8	04-.bwa.drm.sorted.bam|8	3511.45
chr13	28622254	21+0-	chr13	28622305	54+71-	DEL	216	99	67	04-.bwa.drm.sorted.bam|67	3641.50
chr13	28623185	4+0-	chr13	28623267	111+94-	DEL	214	99	89	04-.bwa.drm.sorted.bam|89	188.74
chr13	28624076	111+94-	chr13	28624127	33+25-	DEL	203	99	20	04-.bwa.drm.sorted.bam|20	3338.04
chr13	28624517	33+25-	chr13	28624574	0+5-	DEL	296	99	5	04-.bwa.drm.sorted.bam|5	271.52
chr13	28626641	48+38-	chr13	28627011	48+38-	DEL	228	99	35	04-.bwa.drm.sorted.bam|35	NA
chr13	28631407	7+0-	chr13	28631458	10+14-	DEL	193	99	13	04-.bwa.drm.sorted.bam|13	16386.75
chr13	28631702	10+14-	chr13	28631754	0+2-	DEL	240	79	2	04-.bwa.drm.sorted.bam|2	595.25
chr13	28635911	31+22-	chr13	28636176	31+22-	DEL	190	99	16	04-.bwa.drm.sorted.bam|16	NA
chr13	28636176	31+22-	chr13	28636283	0+3-	DEL	196	99	3	04-.bwa.drm.sorted.bam|3	2024.95
chr13	28644487	71+27-	chr13	28644726	71+27-	DEL	201	99	21	04-.bwa.drm.sorted.bam|21	NA
chr13	28644726	71+27-	chr13	28644783	0+33-	DEL	215	99	33	04-.bwa.drm.sorted.bam|33	8145.46
chr13	28644871	71+27-	chr13	28644931	0+2-	DEL	231	73	2	04-.bwa.drm.sorted.bam|2	7473.96
chr13	28674692	2+0-	chr13	28674708	0+2-	DEL	157	99	2	04-.bwa.drm.sorted.bam|2	2210.91
chr13	29546568	14+5-	chr13	29546710	14+5-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	29546710	14+5-	chr13	29546802	0+8-	DEL	217	99	8	04-.bwa.drm.sorted.bam|8	2523.32
chr13	29546855	14+5-	chr13	29546980	0+3-	DEL	208	99	3	04-.bwa.drm.sorted.bam|3	1433.00
chr13	29735515	2+0-	chr13	29735553	27+25-	DEL	207	99	12	04-.bwa.drm.sorted.bam|12	1183.98
chr13	29735456	7+0-	chr13	29735553	27+25-	DEL	186	99	7	04-.bwa.drm.sorted.bam|7	1116.85
chr13	29735920	27+25-	chr13	29736029	0+2-	DEL	294	73	2	04-.bwa.drm.sorted.bam|2	141.99
chr13	29829047	2+0-	chr13	29829188	41+37-	DEL	204	99	36	04-.bwa.drm.sorted.bam|36	439.05
chr13	30439210	6+0-	chr13	30439244	18+18-	DEL	213	99	12	04-.bwa.drm.sorted.bam|12	2593.81
chr13	30439153	3+0-	chr13	30439244	18+18-	DEL	189	99	3	04-.bwa.drm.sorted.bam|3	3911.61
chr13	31222675	21+11-	chr13	31222791	21+11-	DEL	176	99	6	04-.bwa.drm.sorted.bam|6	NA
chr13	31222791	21+11-	chr13	31222899	0+4-	DEL	201	99	4	04-.bwa.drm.sorted.bam|4	2006.20
chr13	31311958	12+11-	chr13	31312175	12+11-	DEL	186	99	8	04-.bwa.drm.sorted.bam|8	NA
chr13	31596424	15+9-	chr13	31596498	15+9-	DEL	175	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	31950583	6+2-	chr13	31950721	0+3-	DEL	191	99	3	04-.bwa.drm.sorted.bam|3	2467.25
chr13	32242151	13+0-	chr13	32242227	33+32-	DEL	214	99	27	04-.bwa.drm.sorted.bam|27	1018.18
chr13	32242523	33+32-	chr13	32242584	0+10-	DEL	229	99	10	04-.bwa.drm.sorted.bam|10	3805.67
chr13	32390308	10+0-	chr13	32390408	12+15-	DEL	205	99	13	04-.bwa.drm.sorted.bam|13	1083.35
chr13	32773416	13+6-	chr13	32773607	13+6-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	33430809	5+0-	chr13	33430890	8+8-	DEL	199	99	6	04-.bwa.drm.sorted.bam|6	4967.72
chr13	33431084	8+8-	chr13	33431204	0+2-	DEL	174	80	2	04-.bwa.drm.sorted.bam|2	1547.64
chr13	33679831	2+0-	chr13	33679920	23+17-	DEL	203	99	13	04-.bwa.drm.sorted.bam|13	173.89
chr13	33680278	23+17-	chr13	33680372	0+2-	DEL	266	74	2	04-.bwa.drm.sorted.bam|2	658.57
chr13	33691778	35+0-	chr13	33691832	13+44-	DEL	242	99	43	04-.bwa.drm.sorted.bam|43	6018.59
chr13	33787260	3+0-	chr13	33787342	25+22-	DEL	190	99	20	04-.bwa.drm.sorted.bam|20	3208.52
chr13	33946930	31+27-	chr13	33947449	31+27-	DEL	222	99	26	04-.bwa.drm.sorted.bam|26	NA
chr13	34319426	48+36-	chr13	34319782	48+36-	DEL	212	99	32	04-.bwa.drm.sorted.bam|32	NA
chr13	35183178	3+0-	chr13	35183287	17+30-	DEL	218	99	16	04-.bwa.drm.sorted.bam|16	1766.99
chr13	35183226	12+0-	chr13	35183287	17+30-	DEL	199	99	12	04-.bwa.drm.sorted.bam|12	3298.24
chr13	36194227	9+0-	chr13	36194290	6+11-	DEL	204	99	9	04-.bwa.drm.sorted.bam|9	15230.71
chr13	36515140	5+0-	chr13	36515223	6+4-	DEL	187	99	3	04-.bwa.drm.sorted.bam|3	8204.34
chr13	38086939	24+0-	chr13	38086991	15+33-	DEL	221	99	30	04-.bwa.drm.sorted.bam|30	3273.85
chr13	38203403	17+3-	chr13	38203464	17+3-	DEL	174	82	2	04-.bwa.drm.sorted.bam|2	NA
chr13	38203464	17+3-	chr13	38203596	0+2-	DEL	177	81	2	04-.bwa.drm.sorted.bam|2	2931.13
chr13	38730703	12+3-	chr13	38730757	3+11-	DEL	193	99	9	04-.bwa.drm.sorted.bam|9	12610.38
chr13	38730865	3+11-	chr13	38730947	0+2-	DEL	190	88	2	04-.bwa.drm.sorted.bam|2	1321.15
chr13	38733977	11+1-	chr13	38734030	1+10-	DEL	188	99	10	04-.bwa.drm.sorted.bam|10	8176.20
chr13	39000664	8+0-	chr13	39000749	15+15-	DEL	230	99	15	04-.bwa.drm.sorted.bam|15	546.22
chr13	39001046	15+15-	chr13	39001152	0+4-	DEL	232	99	4	04-.bwa.drm.sorted.bam|4	438.01
chr13	39303967	3+0-	chr13	39304094	11+5-	DEL	180	99	3	04-.bwa.drm.sorted.bam|3	1584.20
chr13	39304285	11+5-	chr13	39304380	0+5-	DEL	230	99	5	04-.bwa.drm.sorted.bam|5	814.55
chr13	39304430	11+5-	chr13	39304501	0+3-	DEL	256	99	3	04-.bwa.drm.sorted.bam|3	859.80
chr13	39321238	6+0-	chr13	39321312	5+7-	DEL	191	99	6	04-.bwa.drm.sorted.bam|6	8156.47
chr13	39858204	3+0-	chr13	39858310	12+18-	DEL	250	99	7	04-.bwa.drm.sorted.bam|7	4501.10
chr13	39858239	10+0-	chr13	39858310	12+18-	DEL	193	99	9	04-.bwa.drm.sorted.bam|9	9373.01
chr13	40146143	16+12-	chr13	40146286	16+12-	DEL	181	99	9	04-.bwa.drm.sorted.bam|9	NA
chr13	40146286	16+12-	chr13	40146401	0+3-	DEL	166	99	3	04-.bwa.drm.sorted.bam|3	2018.66
chr13	40432561	16+4-	chr13	40432706	16+4-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	40432706	16+4-	chr13	40432759	0+7-	DEL	188	99	6	04-.bwa.drm.sorted.bam|6	2044.05
chr13	40704597	5+0-	chr13	40704658	12+6-	DEL	182	99	4	04-.bwa.drm.sorted.bam|4	7103.91
chr13	40704824	12+6-	chr13	40704877	0+5-	DEL	174	99	4	04-.bwa.drm.sorted.bam|4	8176.20
chr13	40705535	2+0-	chr13	40705541	28+33-	DEL	212	99	27	04-.bwa.drm.sorted.bam|27	512.46
chr13	40705487	4+0-	chr13	40705541	28+33-	DEL	208	99	4	04-.bwa.drm.sorted.bam|4	286.60
chr13	40786032	10+0-	chr13	40786098	26+12-	DEL	188	99	9	04-.bwa.drm.sorted.bam|9	4455.32
chr13	40786225	26+12-	chr13	40786308	0+15-	DEL	188	99	14	04-.bwa.drm.sorted.bam|14	5780.33
chr13	41196138	4+0-	chr13	41196201	27+22-	DEL	204	99	20	04-.bwa.drm.sorted.bam|20	2210.91
chr13	41215472	2+0-	chr13	41215538	13+9-	DEL	177	99	8	04-.bwa.drm.sorted.bam|8	468.98
chr13	41215776	13+9-	chr13	41215844	0+2-	DEL	215	79	2	04-.bwa.drm.sorted.bam|2	227.59
chr13	41373914	7+0-	chr13	41374014	12+10-	DEL	244	99	8	04-.bwa.drm.sorted.bam|8	2785.75
chr13	41374189	12+10-	chr13	41374251	0+4-	DEL	185	99	4	04-.bwa.drm.sorted.bam|4	7238.95
chr13	42709895	2+0-	chr13	42710014	16+5-	DEL	210	99	3	04-.bwa.drm.sorted.bam|3	520.21
chr13	42710211	16+5-	chr13	42710326	0+11-	DEL	265	99	11	04-.bwa.drm.sorted.bam|11	2287.81
chr13	42782590	5+0-	chr13	42782670	13+8-	DEL	211	99	8	04-.bwa.drm.sorted.bam|8	1934.55
chr13	42782903	13+8-	chr13	42782958	0+5-	DEL	207	99	5	04-.bwa.drm.sorted.bam|5	7034.71
chr13	42949123	4+0-	chr13	42949217	12+5-	DEL	164	99	4	04-.bwa.drm.sorted.bam|4	1975.71
chr13	42949340	12+5-	chr13	42949396	0+6-	DEL	166	99	6	04-.bwa.drm.sorted.bam|6	13265.46
chr13	42949485	12+5-	chr13	42949554	0+2-	DEL	184	86	2	04-.bwa.drm.sorted.bam|2	6653.39
chr13	43117601	29+17-	chr13	43117848	29+17-	DEL	183	99	13	04-.bwa.drm.sorted.bam|13	NA
chr13	43117848	29+17-	chr13	43117906	0+7-	DEL	178	99	7	04-.bwa.drm.sorted.bam|7	2935.17
chr13	43147806	14+0-	chr13	43147868	7+18-	DEL	203	99	14	04-.bwa.drm.sorted.bam|14	5990.85
chr13	43388217	8+3-	chr13	43388343	0+2-	DEL	200	84	2	04-.bwa.drm.sorted.bam|2	12405.66
chr13	43425971	2+0-	chr13	43426095	10+5-	DEL	199	84	2	04-.bwa.drm.sorted.bam|2	748.86
chr13	43426256	10+5-	chr13	43426312	0+3-	DEL	171	99	3	04-.bwa.drm.sorted.bam|3	7185.46
chr13	43944615	8+5-	chr13	43944635	8+5-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	43944780	8+5-	chr13	43944830	0+4-	DEL	204	92	2	04-.bwa.drm.sorted.bam|2	9523.92
chr13	43944736	7+1-	chr13	43944830	0+4-	DEL	173	89	2	04-.bwa.drm.sorted.bam|2	6421.05
chr13	44259726	17+9-	chr13	44259876	17+9-	DEL	193	99	9	04-.bwa.drm.sorted.bam|9	NA
chr13	44259876	17+9-	chr13	44259992	0+2-	DEL	263	75	2	04-.bwa.drm.sorted.bam|2	933.92
chr13	44851864	2+0-	chr13	44851884	17+8-	DEL	212	99	5	04-.bwa.drm.sorted.bam|5	3001.48
chr13	44907447	17+4-	chr13	44907590	17+4-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	44907590	17+4-	chr13	44907695	0+8-	DEL	190	99	8	04-.bwa.drm.sorted.bam|8	3684.85
chr13	44907735	17+4-	chr13	44907825	0+2-	DEL	267	85	2	04-.bwa.drm.sorted.bam|2	2700.13
chr13	45342505	4+0-	chr13	45342602	11+11-	DEL	198	99	10	04-.bwa.drm.sorted.bam|10	1914.60
chr13	45404137	3+0-	chr13	45404260	14+5-	DEL	196	99	3	04-.bwa.drm.sorted.bam|3	880.77
chr13	45404385	14+5-	chr13	45404480	0+6-	DEL	182	99	6	04-.bwa.drm.sorted.bam|6	10426.19
chr13	45404530	14+5-	chr13	45404599	0+4-	DEL	258	99	4	04-.bwa.drm.sorted.bam|4	6870.35
chr13	45997217	12+3-	chr13	45997338	12+3-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	45997338	12+3-	chr13	45997479	0+2-	DEL	184	84	2	04-.bwa.drm.sorted.bam|2	2963.56
chr13	46006214	2+0-	chr13	46006267	20+10-	DEL	184	99	8	04-.bwa.drm.sorted.bam|8	292.01
chr13	46006524	20+10-	chr13	46006582	0+7-	DEL	200	99	7	04-.bwa.drm.sorted.bam|7	2935.17
chr13	46490931	5+0-	chr13	46490982	13+15-	DEL	183	99	13	04-.bwa.drm.sorted.bam|13	10924.50
chr13	46833424	41+37-	chr13	46833876	41+37-	DEL	221	99	35	04-.bwa.drm.sorted.bam|35	NA
chr13	47125530	30+29-	chr13	47125811	30+29-	DEL	201	99	28	04-.bwa.drm.sorted.bam|28	NA
chr13	47236727	2+0-	chr13	47236800	40+5-	DEL	189	99	3	04-.bwa.drm.sorted.bam|3	1060.03
chr13	47236995	40+5-	chr13	47237059	0+27-	DEL	202	99	26	04-.bwa.drm.sorted.bam|26	4110.91
chr13	47706585	18+2-	chr13	47706639	0+16-	DEL	235	99	16	04-.bwa.drm.sorted.bam|16	10030.98
chr13	47837675	26+24-	chr13	47837974	26+24-	DEL	199	99	24	04-.bwa.drm.sorted.bam|24	NA
chr13	48197470	26+3-	chr13	48197543	0+17-	DEL	202	99	16	04-.bwa.drm.sorted.bam|16	9540.23
chr13	49173306	27+19-	chr13	49173522	27+19-	DEL	201	99	17	04-.bwa.drm.sorted.bam|17	NA
chr13	49173522	27+19-	chr13	49173578	0+6-	DEL	239	99	6	04-.bwa.drm.sorted.bam|6	5803.64
chr13	49197434	2+0-	chr13	49197885	14+10-	ITX	-12	99	7	04-.bwa.drm.sorted.bam|7	995.15
chr13	49253401	8+0-	chr13	49253408	4+9-	DEL	179	99	8	04-.bwa.drm.sorted.bam|8	6007.28
chr13	49417847	19+15-	chr13	49418153	19+15-	DEL	198	99	14	04-.bwa.drm.sorted.bam|14	NA
chr13	49434375	3+0-	chr13	49434483	11+4-	DEL	205	99	3	04-.bwa.drm.sorted.bam|3	1576.30
chr13	49434637	11+4-	chr13	49434711	0+5-	DEL	215	99	5	04-.bwa.drm.sorted.bam|5	5228.50
chr13	50098669	2+0-	chr13	50098754	10+9-	DEL	180	99	6	04-.bwa.drm.sorted.bam|6	546.22
chr13	50099108	10+9-	chr13	50099154	0+2-	DEL	217	80	2	04-.bwa.drm.sorted.bam|2	1782.62
chr13	50101093	35+2-	chr13	50101149	0+29-	DEL	209	99	30	04-.bwa.drm.sorted.bam|30	6632.73
chr13	50102610	32+0-	chr13	50102661	8+33-	DEL	211	99	31	04-.bwa.drm.sorted.bam|31	3338.04
chr13	50105760	2+0-	chr13	50105832	39+27-	DEL	213	99	26	04-.bwa.drm.sorted.bam|26	429.90
chr13	50107005	2+0-	chr13	50107135	13+21-	DEL	280	99	3	04-.bwa.drm.sorted.bam|3	5121.27
chr13	50107080	17+0-	chr13	50107135	13+21-	DEL	197	99	17	04-.bwa.drm.sorted.bam|17	14913.59
chr13	50107370	13+21-	chr13	50107435	2+2-	DEL	198	77	2	04-.bwa.drm.sorted.bam|2	476.20
chr13	50107515	13+21-	chr13	50107573	43+36-	DEL	213	99	29	04-.bwa.drm.sorted.bam|29	457.43
chr13	50107497	2+2-	chr13	50107573	43+36-	DEL	310	68	2	04-.bwa.drm.sorted.bam|2	203.64
chr13	50108135	43+36-	chr13	50108191	14+4-	DEL	216	68	2	04-.bwa.drm.sorted.bam|2	6632.73
chr13	50108280	43+36-	chr13	50108337	0+12-	DEL	228	99	5	04-.bwa.drm.sorted.bam|5	10343.12
chr13	50108238	14+4-	chr13	50108337	0+12-	DEL	206	99	7	04-.bwa.drm.sorted.bam|7	6878.39
chr13	51101857	8+0-	chr13	51101920	7+9-	DEL	180	99	7	04-.bwa.drm.sorted.bam|7	13756.77
chr13	51184693	5+0-	chr13	51184772	17+15-	DEL	176	99	12	04-.bwa.drm.sorted.bam|12	3526.26
chr13	51325172	12+4-	chr13	51325235	12+4-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	51325380	12+4-	chr13	51325399	0+4-	DEL	226	99	4	04-.bwa.drm.sorted.bam|4	5662.09
chr13	51357811	3+1-	chr13	51357836	0+2-	DEL	210	96	2	04-.bwa.drm.sorted.bam|2	17661.27
chr13	51365044	17+10-	chr13	51365290	17+10-	ITX	-13	99	5	04-.bwa.drm.sorted.bam|5	NA
chr13	52023464	15+15-	chr13	52023696	15+15-	DEL	204	99	12	04-.bwa.drm.sorted.bam|12	NA
chr13	53271138	2+0-	chr13	53271187	0+2-	DEL	212	99	2	04-.bwa.drm.sorted.bam|2	79.78
chr13	53306219	23+9-	chr13	53306311	23+9-	DEL	165	99	7	04-.bwa.drm.sorted.bam|7	NA
chr13	53306311	23+9-	chr13	53306379	0+7-	DEL	221	99	7	04-.bwa.drm.sorted.bam|7	2731.12
chr13	53306456	23+9-	chr13	53306480	0+2-	DEL	201	78	2	04-.bwa.drm.sorted.bam|2	2289.40
chr13	53447783	2+0-	chr13	53447819	19+18-	DEL	199	99	13	04-.bwa.drm.sorted.bam|13	1539.09
chr13	53447740	3+0-	chr13	53447819	19+18-	DEL	194	99	3	04-.bwa.drm.sorted.bam|3	2742.65
chr13	53639087	19+3-	chr13	53639144	19+3-	DEL	153	82	2	04-.bwa.drm.sorted.bam|2	NA
chr13	53639144	19+3-	chr13	53639248	0+9-	DEL	239	99	9	04-.bwa.drm.sorted.bam|9	2678.60
chr13	53803126	67+64-	chr13	53803475	67+64-	DEL	205	99	59	04-.bwa.drm.sorted.bam|59	NA
chr13	54066757	10+0-	chr13	54066761	13+11-	DEL	217	99	10	04-.bwa.drm.sorted.bam|10	2596.71
chr13	54066919	13+11-	chr13	54066998	0+5-	DEL	197	99	5	04-.bwa.drm.sorted.bam|5	2742.65
chr13	54503124	53+42-	chr13	54503467	53+42-	DEL	204	99	41	04-.bwa.drm.sorted.bam|41	NA
chr13	54503467	53+42-	chr13	54503598	0+2-	DEL	328	70	2	04-.bwa.drm.sorted.bam|2	236.28
chr13	54531090	3+0-	chr13	54531151	18+17-	DEL	180	99	10	04-.bwa.drm.sorted.bam|10	6850.20
chr13	54897742	2+0-	chr13	54897878	51+53-	DEL	227	99	52	04-.bwa.drm.sorted.bam|52	55.08
chr13	55113847	34+19-	chr13	55114170	34+19-	DEL	211	99	16	04-.bwa.drm.sorted.bam|16	NA
chr13	55114170	34+19-	chr13	55114227	0+9-	DEL	265	99	9	04-.bwa.drm.sorted.bam|9	1900.61
chr13	55270310	17+13-	chr13	55270589	17+13-	DEL	212	99	9	04-.bwa.drm.sorted.bam|9	NA
chr13	55818306	25+17-	chr13	55818631	25+17-	DEL	231	99	11	04-.bwa.drm.sorted.bam|11	NA
chr13	55818631	25+17-	chr13	55818691	0+4-	DEL	250	99	4	04-.bwa.drm.sorted.bam|4	2579.40
chr13	56265488	2+0-	chr13	56265593	15+8-	DEL	176	99	3	04-.bwa.drm.sorted.bam|3	5748.37
chr13	56265803	15+8-	chr13	56265898	0+4-	DEL	216	99	4	04-.bwa.drm.sorted.bam|4	1303.27
chr13	56329408	40+32-	chr13	56329845	40+32-	DEL	211	99	30	04-.bwa.drm.sorted.bam|30	NA
chr13	56329845	40+32-	chr13	56329912	0+2-	DEL	358	68	2	04-.bwa.drm.sorted.bam|2	230.99
chr13	57874172	51+47-	chr13	57874707	51+47-	DEL	225	99	47	04-.bwa.drm.sorted.bam|47	NA
chr13	58668490	13+0-	chr13	58668576	11+16-	DEL	205	99	12	04-.bwa.drm.sorted.bam|12	7198.31
chr13	58776262	16+0-	chr13	58776314	10+21-	DEL	199	99	18	04-.bwa.drm.sorted.bam|18	9821.54
chr13	58776520	10+21-	chr13	58776648	0+2-	DEL	229	80	2	04-.bwa.drm.sorted.bam|2	1209.09
chr13	59759959	9+0-	chr13	59760019	9+13-	DEL	162	99	8	04-.bwa.drm.sorted.bam|8	9027.88
chr13	59760151	9+13-	chr13	59760211	0+4-	DEL	152	99	3	04-.bwa.drm.sorted.bam|3	4127.03
chr13	59924829	14+0-	chr13	59924886	26+33-	DEL	234	99	31	04-.bwa.drm.sorted.bam|31	7059.40
chr13	60420033	40+32-	chr13	60420454	40+32-	DEL	206	99	28	04-.bwa.drm.sorted.bam|28	NA
chr13	60420454	40+32-	chr13	60420527	0+4-	DEL	279	99	4	04-.bwa.drm.sorted.bam|4	212.01
chr13	60465169	36+11-	chr13	60465456	36+11-	DEL	214	99	10	04-.bwa.drm.sorted.bam|10	NA
chr13	60465456	36+11-	chr13	60465581	0+18-	DEL	272	99	18	04-.bwa.drm.sorted.bam|18	1733.35
chr13	60672999	23+18-	chr13	60673244	23+18-	DEL	205	99	17	04-.bwa.drm.sorted.bam|17	NA
chr13	60775961	2+0-	chr13	60776025	48+45-	DEL	217	99	41	04-.bwa.drm.sorted.bam|41	241.82
chr13	60849147	5+1-	chr13	60849171	0+3-	DEL	178	99	3	04-.bwa.drm.sorted.bam|3	5311.42
chr13	60918322	20+5-	chr13	60918434	20+5-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	60918434	20+5-	chr13	60918489	0+2-	DEL	160	85	2	04-.bwa.drm.sorted.bam|2	13788.04
chr13	60924706	21+9-	chr13	60924881	21+9-	DEL	176	99	6	04-.bwa.drm.sorted.bam|6	NA
chr13	60924881	21+9-	chr13	60924947	0+2-	DEL	162	75	2	04-.bwa.drm.sorted.bam|2	468.98
chr13	61195386	5+1-	chr13	61195437	6+4-	DEL	177	99	3	04-.bwa.drm.sorted.bam|3	7283.00
chr13	61195696	6+4-	chr13	61195705	0+3-	DEL	234	99	3	04-.bwa.drm.sorted.bam|3	1909.42
chr13	61975084	14+0-	chr13	61975172	42+50-	DEL	218	99	46	04-.bwa.drm.sorted.bam|46	703.47
chr13	61975563	42+50-	chr13	61975642	0+3-	DEL	367	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	62244704	41+31-	chr13	62244941	41+31-	DEL	200	99	25	04-.bwa.drm.sorted.bam|25	NA
chr13	62245086	41+31-	chr13	62245103	0+2-	DEL	283	72	2	04-.bwa.drm.sorted.bam|2	1050.86
chr13	62660128	2+0-	chr13	62660181	7+2-	DEL	174	86	2	04-.bwa.drm.sorted.bam|2	4380.10
chr13	62660467	7+2-	chr13	62660520	0+3-	DEL	312	99	3	04-.bwa.drm.sorted.bam|3	2266.74
chr13	63252123	6+0-	chr13	63252176	26+22-	DEL	192	99	21	04-.bwa.drm.sorted.bam|21	292.01
chr13	63252708	26+22-	chr13	63252710	0+2-	DEL	320	73	2	04-.bwa.drm.sorted.bam|2	105.28
chr13	63277029	30+9-	chr13	63277235	30+9-	DEL	183	99	9	04-.bwa.drm.sorted.bam|9	NA
chr13	63277235	30+9-	chr13	63277289	0+16-	DEL	224	99	16	04-.bwa.drm.sorted.bam|16	1719.60
chr13	63714848	38+2-	chr13	63714905	0+32-	DEL	218	99	33	04-.bwa.drm.sorted.bam|33	2986.67
chr13	64122461	6+0-	chr13	64122542	15+12-	DEL	208	99	7	04-.bwa.drm.sorted.bam|7	2292.80
chr13	64122713	15+12-	chr13	64122772	0+5-	DEL	197	99	5	04-.bwa.drm.sorted.bam|5	2360.80
chr13	64122858	15+12-	chr13	64122872	0+2-	DEL	298	82	2	04-.bwa.drm.sorted.bam|2	1362.70
chr13	64857551	17+0-	chr13	64857632	7+16-	DEL	175	99	14	04-.bwa.drm.sorted.bam|14	4776.66
chr13	64857696	17+0-	chr13	64857802	0+4-	DEL	288	99	3	04-.bwa.drm.sorted.bam|3	10543.66
chr13	64857875	7+16-	chr13	64857934	0+2-	DEL	240	87	2	04-.bwa.drm.sorted.bam|2	1972.48
chr13	64977588	47+37-	chr13	64978038	47+37-	DEL	216	99	34	04-.bwa.drm.sorted.bam|34	NA
chr13	66069459	49+34-	chr13	66069775	49+34-	DEL	228	99	31	04-.bwa.drm.sorted.bam|31	NA
chr13	66069775	49+34-	chr13	66069838	0+12-	DEL	245	99	12	04-.bwa.drm.sorted.bam|12	2702.22
chr13	66648497	8+0-	chr13	66648637	33+37-	DEL	200	99	31	04-.bwa.drm.sorted.bam|31	1216.00
chr13	66648586	3+0-	chr13	66648637	33+37-	DEL	244	99	3	04-.bwa.drm.sorted.bam|3	1213.83
chr13	66649031	33+37-	chr13	66649105	0+3-	DEL	369	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	67179788	14+0-	chr13	67179893	12+20-	DEL	192	99	19	04-.bwa.drm.sorted.bam|19	1768.73
chr13	67300877	26+0-	chr13	67300934	10+32-	DEL	202	99	31	04-.bwa.drm.sorted.bam|31	12218.19
chr13	67774367	2+0-	chr13	67774395	6+3-	DEL	187	88	2	04-.bwa.drm.sorted.bam|2	984.05
chr13	67904945	3+0-	chr13	67905040	22+12-	DEL	185	99	9	04-.bwa.drm.sorted.bam|9	1629.09
chr13	67905315	22+12-	chr13	67905397	0+7-	DEL	223	99	7	04-.bwa.drm.sorted.bam|7	754.95
chr13	67929906	16+0-	chr13	67929957	12+19-	DEL	171	99	15	04-.bwa.drm.sorted.bam|15	6069.17
chr13	67930243	12+19-	chr13	67930259	0+3-	DEL	199	99	3	04-.bwa.drm.sorted.bam|3	1249.64
chr13	68405821	40+17-	chr13	68406016	40+17-	DEL	200	99	14	04-.bwa.drm.sorted.bam|14	NA
chr13	68406016	40+17-	chr13	68406080	0+15-	DEL	242	99	15	04-.bwa.drm.sorted.bam|15	6529.09
chr13	68948987	2+0-	chr13	68949047	24+22-	DEL	206	99	21	04-.bwa.drm.sorted.bam|21	515.88
chr13	69558981	2+3-	chr13	69559044	2+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	70123493	22+20-	chr13	70123767	22+20-	DEL	203	99	18	04-.bwa.drm.sorted.bam|18	NA
chr13	70265113	27+19-	chr13	70265447	27+19-	DEL	192	99	13	04-.bwa.drm.sorted.bam|13	NA
chr13	70265447	27+19-	chr13	70265580	0+2-	DEL	342	70	2	04-.bwa.drm.sorted.bam|2	116.36
chr13	70286169	29+0-	chr13	70286224	23+35-	DEL	235	99	31	04-.bwa.drm.sorted.bam|31	2251.11
chr13	70286474	23+35-	chr13	70286530	0+12-	DEL	205	99	11	04-.bwa.drm.sorted.bam|11	1658.18
chr13	71118187	24+20-	chr13	71118530	24+20-	DEL	195	99	18	04-.bwa.drm.sorted.bam|18	NA
chr13	71327908	33+32-	chr13	71328331	33+32-	DEL	223	99	30	04-.bwa.drm.sorted.bam|30	NA
chr13	71850931	2+0-	chr13	71850946	6+4-	DEL	228	86	2	04-.bwa.drm.sorted.bam|2	1257.46
chr13	72306070	24+18-	chr13	72306308	24+18-	DEL	191	99	17	04-.bwa.drm.sorted.bam|17	NA
chr13	72306308	24+18-	chr13	72306364	0+3-	DEL	209	99	3	04-.bwa.drm.sorted.bam|3	2487.27
chr13	72332509	12+0-	chr13	72332566	24+27-	DEL	191	99	24	04-.bwa.drm.sorted.bam|24	4344.24
chr13	72341658	35+33-	chr13	72342034	35+33-	DEL	214	99	26	04-.bwa.drm.sorted.bam|26	NA
chr13	72425237	69+60-	chr13	72425690	69+60-	DEL	204	99	59	04-.bwa.drm.sorted.bam|59	NA
chr13	72425690	69+60-	chr13	72425748	17+14-	DEL	194	99	13	04-.bwa.drm.sorted.bam|13	800.50
chr13	73952490	10+4-	chr13	73952553	10+4-	DEL	155	82	2	04-.bwa.drm.sorted.bam|2	NA
chr13	73952553	10+4-	chr13	73952619	0+2-	DEL	184	81	2	04-.bwa.drm.sorted.bam|2	2813.89
chr13	73952553	10+4-	chr13	73952680	0+4-	DEL	187	99	4	04-.bwa.drm.sorted.bam|4	2071.64
chr13	74099765	10+0-	chr13	74099832	11+17-	DEL	194	99	13	04-.bwa.drm.sorted.bam|13	3926.84
chr13	74238074	19+17-	chr13	74238320	19+17-	DEL	187	99	14	04-.bwa.drm.sorted.bam|14	NA
chr13	74336701	12+1-	chr13	74336754	1+10-	DEL	203	99	11	04-.bwa.drm.sorted.bam|11	8176.20
chr13	74373644	16+12-	chr13	74373869	16+12-	DEL	201	99	11	04-.bwa.drm.sorted.bam|11	NA
chr13	74373869	16+12-	chr13	74373958	0+4-	DEL	252	99	4	04-.bwa.drm.sorted.bam|4	1043.35
chr13	74387897	14+0-	chr13	74387958	14+19-	DEL	208	99	15	04-.bwa.drm.sorted.bam|15	10402.15
chr13	74388136	14+19-	chr13	74388196	0+3-	DEL	205	99	3	04-.bwa.drm.sorted.bam|3	3869.09
chr13	74388281	14+19-	chr13	74388336	0+2-	DEL	248	81	2	04-.bwa.drm.sorted.bam|2	1702.40
chr13	74863091	8+0-	chr13	74863165	20+15-	DEL	183	99	12	04-.bwa.drm.sorted.bam|12	2300.54
chr13	74863370	20+15-	chr13	74863500	0+2-	DEL	198	79	2	04-.bwa.drm.sorted.bam|2	1547.64
chr13	75026530	7+0-	chr13	75026595	8+10-	DEL	178	99	7	04-.bwa.drm.sorted.bam|7	21666.92
chr13	75137835	3+0-	chr13	75137906	42+37-	DEL	214	99	34	04-.bwa.drm.sorted.bam|34	217.98
chr13	75138278	42+37-	chr13	75138338	0+2-	DEL	251	74	2	04-.bwa.drm.sorted.bam|2	1031.76
chr13	75681441	2+0-	chr13	75681495	64+62-	DEL	230	99	57	04-.bwa.drm.sorted.bam|57	NA
chr13	75827434	5+3-	chr13	75827527	5+3-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	75827434	5+3-	chr13	75827774	5+5-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	1684.19
chr13	75870467	45+38-	chr13	75870979	45+38-	DEL	231	99	34	04-.bwa.drm.sorted.bam|34	NA
chr13	75870979	45+38-	chr13	75871058	0+3-	DEL	370	91	3	04-.bwa.drm.sorted.bam|3	NA
chr13	75880569	11+7-	chr13	75880645	11+7-	DEL	175	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	75880645	11+7-	chr13	75880703	0+2-	DEL	198	80	2	04-.bwa.drm.sorted.bam|2	2935.17
chr13	75880645	11+7-	chr13	75880774	11+4-	DEL	271	99	4	04-.bwa.drm.sorted.bam|4	1679.61
chr13	75880923	11+4-	chr13	75880992	5+11-	DEL	188	99	10	04-.bwa.drm.sorted.bam|10	15027.78
chr13	76416767	5+0-	chr13	76416897	20+20-	DEL	244	99	16	04-.bwa.drm.sorted.bam|16	1428.59
chr13	76416846	3+0-	chr13	76416897	20+20-	DEL	237	99	3	04-.bwa.drm.sorted.bam|3	2124.21
chr13	76512661	37+31-	chr13	76513043	37+31-	DEL	191	99	27	04-.bwa.drm.sorted.bam|27	NA
chr13	76923209	10+1-	chr13	76923282	4+8-	DEL	200	99	8	04-.bwa.drm.sorted.bam|8	5088.12
chr13	77397921	4+0-	chr13	77397972	9+10-	DEL	173	99	4	04-.bwa.drm.sorted.bam|4	10621.04
chr13	77443488	5+0-	chr13	77443604	4+8-	DEL	174	99	5	04-.bwa.drm.sorted.bam|5	4002.51
chr13	77914802	12+1-	chr13	77914854	2+7-	DEL	166	99	4	04-.bwa.drm.sorted.bam|4	10416.79
chr13	77914947	12+1-	chr13	77914999	0+2-	DEL	233	89	2	04-.bwa.drm.sorted.bam|2	9034.43
chr13	77919643	26+21-	chr13	77919922	26+21-	DEL	199	99	17	04-.bwa.drm.sorted.bam|17	NA
chr13	78023271	2+0-	chr13	78023329	27+8-	DEL	189	99	5	04-.bwa.drm.sorted.bam|5	533.67
chr13	78023558	27+8-	chr13	78023615	0+13-	DEL	222	99	13	04-.bwa.drm.sorted.bam|13	2172.12
chr13	78371661	6+0-	chr13	78371727	18+6-	DEL	169	99	6	04-.bwa.drm.sorted.bam|6	2579.40
chr13	78371861	18+6-	chr13	78371983	0+8-	DEL	215	99	8	04-.bwa.drm.sorted.bam|8	3932.52
chr13	78377599	18+0-	chr13	78377667	21+19-	DEL	199	99	14	04-.bwa.drm.sorted.bam|14	1365.56
chr13	78377744	18+0-	chr13	78377885	0+16-	DEL	372	99	4	04-.bwa.drm.sorted.bam|4	12337.81
chr13	78377830	21+19-	chr13	78377885	0+16-	DEL	203	99	12	04-.bwa.drm.sorted.bam|12	6190.55
chr13	78808915	25+1-	chr13	78809019	0+19-	DEL	231	99	19	04-.bwa.drm.sorted.bam|19	8035.81
chr13	78972506	14+9-	chr13	78972743	14+9-	DEL	210	99	7	04-.bwa.drm.sorted.bam|7	NA
chr13	79172540	27+0-	chr13	79172608	2+27-	DEL	224	99	27	04-.bwa.drm.sorted.bam|27	4324.28
chr13	79699390	8+3-	chr13	79699489	0+5-	DEL	202	99	5	04-.bwa.drm.sorted.bam|5	3439.19
chr13	79920861	67+64-	chr13	79921295	67+64-	DEL	225	99	57	04-.bwa.drm.sorted.bam|57	NA
chr13	80168921	39+2-	chr13	80168987	0+34-	DEL	230	99	34	04-.bwa.drm.sorted.bam|34	19931.69
chr13	81183724	26+17-	chr13	81183937	26+17-	DEL	201	99	11	04-.bwa.drm.sorted.bam|11	NA
chr13	81184082	26+17-	chr13	81184175	0+2-	DEL	284	74	2	04-.bwa.drm.sorted.bam|2	2340.96
chr13	82132468	2+0-	chr13	82132548	11+10-	DEL	208	99	5	04-.bwa.drm.sorted.bam|5	580.36
chr13	82132813	11+10-	chr13	82132891	0+2-	DEL	234	77	2	04-.bwa.drm.sorted.bam|2	1587.32
chr13	84147628	2+0-	chr13	84147708	30+42-	DEL	219	99	26	04-.bwa.drm.sorted.bam|26	1169.33
chr13	84147653	14+0-	chr13	84147708	30+42-	DEL	193	99	14	04-.bwa.drm.sorted.bam|14	562.78
chr13	85202627	28+19-	chr13	85202789	28+19-	DEL	174	99	14	04-.bwa.drm.sorted.bam|14	NA
chr13	85202789	28+19-	chr13	85202896	0+8-	DEL	231	99	8	04-.bwa.drm.sorted.bam|8	3471.34
chr13	85475122	2+0-	chr13	85475230	20+7-	DEL	279	85	2	04-.bwa.drm.sorted.bam|2	1529.29
chr13	85475210	2+0-	chr13	85475230	20+7-	DEL	238	84	2	04-.bwa.drm.sorted.bam|2	2157.31
chr13	85475171	2+0-	chr13	85475230	20+7-	DEL	196	83	2	04-.bwa.drm.sorted.bam|2	4721.60
chr13	85475379	20+7-	chr13	85475498	0+12-	DEL	225	99	12	04-.bwa.drm.sorted.bam|12	4421.82
chr13	86316592	10+0-	chr13	86316649	17+14-	DEL	224	99	12	04-.bwa.drm.sorted.bam|12	271.52
chr13	86316871	17+14-	chr13	86316925	0+10-	DEL	211	99	9	04-.bwa.drm.sorted.bam|9	3439.19
chr13	86317016	17+14-	chr13	86317097	0+3-	DEL	271	99	3	04-.bwa.drm.sorted.bam|3	3218.54
chr13	86740570	20+2-	chr13	86740672	0+10-	DEL	191	99	10	04-.bwa.drm.sorted.bam|10	15779.83
chr13	86949158	2+0-	chr13	86949230	47+49-	DEL	222	99	44	04-.bwa.drm.sorted.bam|44	214.95
chr13	88545286	2+0-	chr13	88545383	19+18-	DEL	223	99	4	04-.bwa.drm.sorted.bam|4	2877.84
chr13	88545317	12+0-	chr13	88545383	19+18-	DEL	189	99	11	04-.bwa.drm.sorted.bam|11	4924.30
chr13	88545706	19+18-	chr13	88545763	0+2-	DEL	260	83	2	04-.bwa.drm.sorted.bam|2	1302.47
chr13	89229851	6+0-	chr13	89229930	22+21-	DEL	209	99	17	04-.bwa.drm.sorted.bam|17	195.90
chr13	89636843	45+29-	chr13	89637099	45+29-	DEL	217	99	24	04-.bwa.drm.sorted.bam|24	NA
chr13	89637099	45+29-	chr13	89637157	0+10-	DEL	236	99	10	04-.bwa.drm.sorted.bam|10	1334.17
chr13	89637244	45+29-	chr13	89637314	0+2-	DEL	325	72	2	04-.bwa.drm.sorted.bam|2	1151.73
chr13	90338888	14+8-	chr13	90339033	14+8-	DEL	182	99	7	04-.bwa.drm.sorted.bam|7	NA
chr13	90822867	28+24-	chr13	90823091	28+24-	DEL	189	99	17	04-.bwa.drm.sorted.bam|17	NA
chr13	91152985	27+14-	chr13	91153230	27+14-	DEL	192	99	12	04-.bwa.drm.sorted.bam|12	NA
chr13	91153230	27+14-	chr13	91153297	0+3-	DEL	248	99	3	04-.bwa.drm.sorted.bam|3	923.96
chr13	92015716	42+33-	chr13	92016137	42+33-	DEL	220	99	29	04-.bwa.drm.sorted.bam|29	NA
chr13	92016137	42+33-	chr13	92016194	0+4-	DEL	328	99	4	04-.bwa.drm.sorted.bam|4	271.52
chr13	92107985	4+0-	chr13	92108096	16+9-	DEL	173	99	4	04-.bwa.drm.sorted.bam|4	3067.39
chr13	92108200	16+9-	chr13	92108264	0+7-	DEL	213	99	6	04-.bwa.drm.sorted.bam|6	14509.10
chr13	92121260	26+8-	chr13	92121379	26+8-	DEL	181	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	92121379	26+8-	chr13	92121448	0+4-	DEL	182	99	4	04-.bwa.drm.sorted.bam|4	1570.07
chr13	92122302	30+16-	chr13	92122530	30+16-	DEL	193	99	15	04-.bwa.drm.sorted.bam|15	NA
chr13	92122530	30+16-	chr13	92122584	0+11-	DEL	257	99	11	04-.bwa.drm.sorted.bam|11	3152.59
chr13	92137196	11+2-	chr13	92137312	11+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	92137312	11+2-	chr13	92137452	0+4-	DEL	177	99	4	04-.bwa.drm.sorted.bam|4	5306.18
chr13	92140223	3+0-	chr13	92140344	10+5-	DEL	164	99	3	04-.bwa.drm.sorted.bam|3	2941.79
chr13	92140410	10+5-	chr13	92140467	1+8-	DEL	183	99	7	04-.bwa.drm.sorted.bam|7	15204.86
chr13	92142118	3+0-	chr13	92142193	9+6-	DEL	182	99	3	04-.bwa.drm.sorted.bam|3	7222.31
chr13	92142459	9+6-	chr13	92142521	0+3-	DEL	262	99	3	04-.bwa.drm.sorted.bam|3	822.42
chr13	92239073	19+0-	chr13	92239124	21+21-	DEL	221	99	19	04-.bwa.drm.sorted.bam|19	3034.58
chr13	92239322	21+21-	chr13	92239374	0+10-	DEL	199	99	9	04-.bwa.drm.sorted.bam|9	3273.85
chr13	92260109	32+0-	chr13	92260176	16+31-	DEL	195	99	27	04-.bwa.drm.sorted.bam|27	6005.76
chr13	92260254	32+0-	chr13	92260356	0+8-	DEL	307	99	5	04-.bwa.drm.sorted.bam|5	16478.89
chr13	92260300	16+31-	chr13	92260356	0+8-	DEL	175	99	3	04-.bwa.drm.sorted.bam|3	8290.91
chr13	92379319	3+0-	chr13	92379438	24+11-	DEL	197	99	10	04-.bwa.drm.sorted.bam|10	3771.55
chr13	92379694	24+11-	chr13	92379749	0+9-	DEL	215	99	9	04-.bwa.drm.sorted.bam|9	844.17
chr13	92379839	24+11-	chr13	92379889	0+3-	DEL	336	99	3	04-.bwa.drm.sorted.bam|3	952.39
chr13	92732695	11+0-	chr13	92732746	25+24-	DEL	246	99	17	04-.bwa.drm.sorted.bam|17	910.37
chr13	92733008	25+24-	chr13	92733077	0+4-	DEL	192	99	4	04-.bwa.drm.sorted.bam|4	2018.66
chr13	92733153	25+24-	chr13	92733274	0+2-	DEL	392	77	2	04-.bwa.drm.sorted.bam|2	930.91
chr13	92891273	10+0-	chr13	92891331	55+65-	DEL	205	99	62	04-.bwa.drm.sorted.bam|62	1067.34
chr13	92892097	30+24-	chr13	92892372	30+24-	DEL	194	99	23	04-.bwa.drm.sorted.bam|23	NA
chr13	92892372	30+24-	chr13	92892430	0+3-	DEL	288	99	3	04-.bwa.drm.sorted.bam|3	533.67
chr13	92902238	21+15-	chr13	92902396	21+15-	DEL	185	99	12	04-.bwa.drm.sorted.bam|12	NA
chr13	92902396	21+15-	chr13	92902465	0+3-	DEL	247	99	3	04-.bwa.drm.sorted.bam|3	2242.95
chr13	92962502	5+0-	chr13	92962590	16+6-	DEL	210	99	3	04-.bwa.drm.sorted.bam|3	4220.83
chr13	92962647	5+0-	chr13	92962800	0+8-	DEL	334	85	2	04-.bwa.drm.sorted.bam|2	11425.51
chr13	92962740	16+6-	chr13	92962800	0+8-	DEL	203	99	6	04-.bwa.drm.sorted.bam|6	3869.09
chr13	92970710	5+1-	chr13	92970725	0+4-	DEL	221	99	4	04-.bwa.drm.sorted.bam|4	483.64
chr13	92978101	2+0-	chr13	92978193	32+28-	DEL	211	99	27	04-.bwa.drm.sorted.bam|27	168.22
chr13	93279016	43+41-	chr13	93279500	43+41-	DEL	238	99	38	04-.bwa.drm.sorted.bam|38	NA
chr13	93842150	8+0-	chr13	93842202	12+17-	DEL	193	99	14	04-.bwa.drm.sorted.bam|14	3273.85
chr13	94017970	29+26-	chr13	94018303	29+26-	DEL	200	99	24	04-.bwa.drm.sorted.bam|24	NA
chr13	94299379	39+31-	chr13	94299715	39+31-	DEL	201	99	29	04-.bwa.drm.sorted.bam|29	NA
chr13	95147584	33+34-	chr13	95147936	33+34-	DEL	224	99	33	04-.bwa.drm.sorted.bam|33	NA
chr13	95675763	5+0-	chr13	95675872	14+11-	DEL	221	99	5	04-.bwa.drm.sorted.bam|5	8661.09
chr13	95676057	14+11-	chr13	95676145	4+4-	DEL	202	99	4	04-.bwa.drm.sorted.bam|4	3341.49
chr13	95676265	4+4-	chr13	95676335	7+6-	DEL	190	99	6	04-.bwa.drm.sorted.bam|6	884.36
chr13	95676543	7+6-	chr13	95676595	0+4-	DEL	216	99	4	04-.bwa.drm.sorted.bam|4	1190.49
chr13	95731466	3+0-	chr13	95731502	1+3-	DEL	192	99	3	04-.bwa.drm.sorted.bam|3	6327.36
chr13	95731643	21+5-	chr13	95731807	21+5-	ITX	-13	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	95731807	21+5-	chr13	95731882	0+7-	DEL	202	99	7	04-.bwa.drm.sorted.bam|7	2476.22
chr13	95747981	26+6-	chr13	95748115	26+6-	DEL	195	99	5	04-.bwa.drm.sorted.bam|5	NA
chr13	95748115	26+6-	chr13	95748175	6+20-	DEL	261	99	19	04-.bwa.drm.sorted.bam|19	12896.98
chr13	95748319	6+20-	chr13	95748437	0+3-	DEL	195	99	3	04-.bwa.drm.sorted.bam|3	262.31
chr13	95785511	3+0-	chr13	95785573	10+11-	DEL	201	99	6	04-.bwa.drm.sorted.bam|6	9735.14
chr13	96159289	13+0-	chr13	96159423	7+15-	DEL	188	99	11	04-.bwa.drm.sorted.bam|11	2309.91
chr13	96159434	13+0-	chr13	96159585	0+4-	DEL	311	86	2	04-.bwa.drm.sorted.bam|2	6378.77
chr13	96159524	7+15-	chr13	96159666	0+4-	DEL	171	99	4	04-.bwa.drm.sorted.bam|4	5340.44
chr13	97040316	10+0-	chr13	97040376	13+10-	DEL	195	99	9	04-.bwa.drm.sorted.bam|9	5416.73
chr13	97040530	13+10-	chr13	97040585	0+3-	DEL	185	82	2	04-.bwa.drm.sorted.bam|2	3939.44
chr13	97465338	22+20-	chr13	97465584	22+20-	DEL	205	99	18	04-.bwa.drm.sorted.bam|18	NA
chr13	98244176	8+6-	chr13	98244307	8+6-	ITX	-10	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	98314257	20+16-	chr13	98314475	20+16-	DEL	184	99	10	04-.bwa.drm.sorted.bam|10	NA
chr13	99398713	34+23-	chr13	99398989	34+23-	DEL	200	99	22	04-.bwa.drm.sorted.bam|22	NA
chr13	99398989	34+23-	chr13	99399044	0+4-	DEL	222	99	4	04-.bwa.drm.sorted.bam|4	2813.89
chr13	99401492	2+0-	chr13	99401583	31+8-	DEL	220	99	6	04-.bwa.drm.sorted.bam|6	170.07
chr13	99401851	31+8-	chr13	99401981	0+13-	DEL	208	99	13	04-.bwa.drm.sorted.bam|13	2500.03
chr13	100645525	7+0-	chr13	100645546	20+17-	DEL	262	99	9	04-.bwa.drm.sorted.bam|9	2144.32
chr13	100645474	8+0-	chr13	100645546	20+17-	DEL	223	99	7	04-.bwa.drm.sorted.bam|7	1719.60
chr13	100645746	20+17-	chr13	100645862	0+9-	DEL	182	99	8	04-.bwa.drm.sorted.bam|8	3202.01
chr13	100645891	20+17-	chr13	100646018	0+4-	DEL	331	99	4	04-.bwa.drm.sorted.bam|4	1820.75
chr13	100895770	3+0-	chr13	100895850	2+4-	DEL	164	88	2	04-.bwa.drm.sorted.bam|2	4256.00
chr13	101571854	4+0-	chr13	101571892	27+23-	DEL	222	99	14	04-.bwa.drm.sorted.bam|14	845.70
chr13	101571820	4+0-	chr13	101571892	27+23-	DEL	207	99	4	04-.bwa.drm.sorted.bam|4	1074.75
chr13	101572135	27+23-	chr13	101572217	0+5-	DEL	231	99	5	04-.bwa.drm.sorted.bam|5	566.21
chr13	101723791	30+25-	chr13	101724216	30+25-	DEL	195	99	21	04-.bwa.drm.sorted.bam|21	NA
chr13	101795230	40+37-	chr13	101795587	40+37-	DEL	201	99	33	04-.bwa.drm.sorted.bam|33	NA
chr13	102518456	37+0-	chr13	102518535	7+36-	DEL	262	99	35	04-.bwa.drm.sorted.bam|35	3134.45
chr13	102518601	37+0-	chr13	102518720	0+4-	DEL	283	75	2	04-.bwa.drm.sorted.bam|2	14890.14
chr13	102518662	7+36-	chr13	102518720	0+4-	DEL	192	86	2	04-.bwa.drm.sorted.bam|2	5069.85
chr13	102696069	14+8-	chr13	102696279	14+8-	ITX	-12	99	5	04-.bwa.drm.sorted.bam|5	NA
chr13	102696279	14+8-	chr13	102696367	0+2-	DEL	172	80	2	04-.bwa.drm.sorted.bam|2	2813.89
chr13	103350468	2+0-	chr13	103350560	8+5-	DEL	177	99	4	04-.bwa.drm.sorted.bam|4	2355.10
chr13	103350797	8+5-	chr13	103350872	0+2-	DEL	162	79	2	04-.bwa.drm.sorted.bam|2	3095.27
chr13	103504085	2+0-	chr13	103504168	56+50-	DEL	239	99	49	04-.bwa.drm.sorted.bam|49	67.88
chr13	103504842	56+50-	chr13	103504925	0+2-	DEL	380	66	2	04-.bwa.drm.sorted.bam|2	186.46
chr13	103683174	8+0-	chr13	103683231	15+15-	DEL	208	99	14	04-.bwa.drm.sorted.bam|14	1086.06
chr13	103683498	15+15-	chr13	103683562	0+3-	DEL	209	99	3	04-.bwa.drm.sorted.bam|3	3627.27
chr13	103684867	26+17-	chr13	103685197	26+17-	DEL	199	99	16	04-.bwa.drm.sorted.bam|16	NA
chr13	103914098	12+0-	chr13	103914170	13+12-	DEL	230	99	11	04-.bwa.drm.sorted.bam|11	2149.50
chr13	103914309	13+12-	chr13	103914372	4+11-	DEL	184	99	8	04-.bwa.drm.sorted.bam|8	5404.45
chr13	103914605	4+11-	chr13	103914606	0+2-	DEL	222	90	2	04-.bwa.drm.sorted.bam|2	212.01
chr13	104490683	14+10-	chr13	104490832	14+10-	DEL	195	99	6	04-.bwa.drm.sorted.bam|6	NA
chr13	104490832	14+10-	chr13	104490908	0+3-	DEL	200	99	3	04-.bwa.drm.sorted.bam|3	203.64
chr13	104492346	39+32-	chr13	104492723	39+32-	DEL	230	99	30	04-.bwa.drm.sorted.bam|30	NA
chr13	104665106	33+19-	chr13	104665371	33+19-	DEL	194	99	18	04-.bwa.drm.sorted.bam|18	NA
chr13	104665371	33+19-	chr13	104665428	0+12-	DEL	288	99	12	04-.bwa.drm.sorted.bam|12	1086.06
chr13	104951521	14+0-	chr13	104951648	13+17-	DEL	206	99	14	04-.bwa.drm.sorted.bam|14	4265.14
chr13	104951818	13+17-	chr13	104951875	0+8-	DEL	193	99	8	04-.bwa.drm.sorted.bam|8	2986.67
chr13	105464629	37+0-	chr13	105464692	5+37-	DEL	223	99	36	04-.bwa.drm.sorted.bam|36	3439.19
chr13	105555788	33+29-	chr13	105556338	33+29-	DEL	224	99	28	04-.bwa.drm.sorted.bam|28	NA
chr13	105864099	2+0-	chr13	105864502	10+5-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	921.67
chr13	106032599	2+0-	chr13	106032655	43+38-	DEL	194	99	38	04-.bwa.drm.sorted.bam|38	276.36
chr13	106386434	3+1-	chr13	106386503	4+4-	DEL	159	90	2	04-.bwa.drm.sorted.bam|2	6728.86
chr13	106632341	36+9-	chr13	106632495	36+9-	DEL	189	99	8	04-.bwa.drm.sorted.bam|8	NA
chr13	106632495	36+9-	chr13	106632553	0+27-	DEL	278	99	27	04-.bwa.drm.sorted.bam|27	1867.84
chr13	106651451	17+12-	chr13	106651655	17+12-	DEL	197	99	10	04-.bwa.drm.sorted.bam|10	NA
chr13	106843867	34+23-	chr13	106844213	34+23-	DEL	228	99	21	04-.bwa.drm.sorted.bam|21	NA
chr13	106844358	34+23-	chr13	106844374	0+6-	DEL	235	99	6	04-.bwa.drm.sorted.bam|6	961.27
chr13	107014007	6+0-	chr13	107014065	56+62-	DEL	202	99	57	04-.bwa.drm.sorted.bam|57	800.50
chr13	107579319	19+6-	chr13	107579481	19+6-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	NA
chr13	107579481	19+6-	chr13	107579609	0+4-	DEL	184	99	4	04-.bwa.drm.sorted.bam|4	2660.00
chr13	108612517	12+0-	chr13	108612580	18+14-	DEL	191	99	12	04-.bwa.drm.sorted.bam|12	7369.70
chr13	108612709	18+14-	chr13	108612822	0+4-	DEL	204	99	4	04-.bwa.drm.sorted.bam|4	3013.10
chr13	108668168	2+0-	chr13	108668394	9+19-	DEL	334	99	3	04-.bwa.drm.sorted.bam|3	3253.79
chr13	108668273	7+0-	chr13	108668394	9+19-	DEL	294	99	7	04-.bwa.drm.sorted.bam|7	4130.91
chr13	108668313	9+0-	chr13	108668394	9+19-	DEL	226	99	8	04-.bwa.drm.sorted.bam|8	10508.65
chr13	108668605	9+19-	chr13	108668683	0+4-	DEL	199	99	3	04-.bwa.drm.sorted.bam|3	992.08
chr13	109069025	43+40-	chr13	109069495	43+40-	DEL	214	99	39	04-.bwa.drm.sorted.bam|39	NA
chr13	109374381	5+0-	chr13	109374496	28+32-	DEL	218	99	20	04-.bwa.drm.sorted.bam|20	2826.12
chr13	109374445	4+0-	chr13	109374496	28+32-	DEL	194	99	4	04-.bwa.drm.sorted.bam|4	4248.42
chr13	109703749	44+42-	chr13	109704185	44+42-	DEL	211	99	39	04-.bwa.drm.sorted.bam|39	NA
chr13	109727909	36+24-	chr13	109728187	36+24-	DEL	197	99	18	04-.bwa.drm.sorted.bam|18	NA
chr13	109728187	36+24-	chr13	109728240	0+5-	DEL	314	99	5	04-.bwa.drm.sorted.bam|5	876.02
chr13	109747619	14+2-	chr13	109747716	14+2-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	109747716	14+2-	chr13	109747834	0+3-	DEL	195	99	3	04-.bwa.drm.sorted.bam|3	3803.52
chr13	110823321	14+8-	chr13	110823430	14+8-	DEL	185	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	110936078	14+3-	chr13	110936187	14+3-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	110936187	14+3-	chr13	110936253	0+3-	DEL	174	84	2	04-.bwa.drm.sorted.bam|2	8910.64
chr13	111081980	21+17-	chr13	111082193	21+17-	DEL	207	99	13	04-.bwa.drm.sorted.bam|13	NA
chr13	111117508	13+3-	chr13	111117697	13+3-	ITX	-14	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	111117697	13+3-	chr13	111117767	0+8-	DEL	188	99	8	04-.bwa.drm.sorted.bam|8	5748.37
chr13	111467505	33+31-	chr13	111467913	33+31-	DEL	210	99	30	04-.bwa.drm.sorted.bam|30	NA
chr13	111575606	2+0-	chr13	111575732	12+9-	DEL	205	99	8	04-.bwa.drm.sorted.bam|8	1473.94
chr13	111668513	3+0-	chr13	111668568	5+5-	DEL	201	99	3	04-.bwa.drm.sorted.bam|3	15757.76
chr13	111686142	3+2-	chr13	111686156	3+2-	ITX	-10	99	2	04-.bwa.drm.sorted.bam|2	NA
chr13	112225059	45+36-	chr13	112225349	45+36-	DEL	190	99	35	04-.bwa.drm.sorted.bam|35	NA
chr13	112570252	25+5-	chr13	112570348	25+5-	DEL	174	99	3	04-.bwa.drm.sorted.bam|3	NA
chr13	112570348	25+5-	chr13	112570399	0+11-	DEL	213	99	11	04-.bwa.drm.sorted.bam|11	6069.17
chr13	113293417	11+3-	chr13	113293503	11+3-	DEL	168	80	2	04-.bwa.drm.sorted.bam|2	NA
chr13	113293503	11+3-	chr13	113293601	0+2-	DEL	217	79	2	04-.bwa.drm.sorted.bam|2	5527.28
chr13	113674386	9+0-	chr13	113674457	5+11-	DEL	164	99	8	04-.bwa.drm.sorted.bam|8	19835.91
chr13	114527639	7+0-	chr13	114527713	10+16-	DEL	191	99	11	04-.bwa.drm.sorted.bam|11	16522.07
chr13	114527927	10+16-	chr13	114528045	0+2-	DEL	206	79	2	04-.bwa.drm.sorted.bam|2	131.16
chr13	114843532	2+0-	chr13	114843639	15+4-	DEL	195	85	2	04-.bwa.drm.sorted.bam|2	1880.31
chr13	114843768	15+4-	chr13	114843825	0+3-	DEL	195	99	3	04-.bwa.drm.sorted.bam|3	10317.58
chr13	114843913	15+4-	chr13	114843951	0+6-	DEL	208	99	6	04-.bwa.drm.sorted.bam|6	5919.92
chr14	23586792	3+0-	chr14	23586905	0+2-	DEL	184	98	2	04-.bwa.drm.sorted.bam|2	4858.86
chr14	96854202	3+0-	chr14	96854216	0+2-	DEL	178	98	2	04-.bwa.drm.sorted.bam|2	681.35
chr14	102309367	2+0-	chr14	102309418	32+31-	DEL	229	99	25	04-.bwa.drm.sorted.bam|25	303.46
chr14	102702012	2+0-	chr14	102702140	2+4-	DEL	294	92	2	04-.bwa.drm.sorted.bam|2	1814.08
chr15	20945754	40+22-	chr15	20945974	40+22-	DEL	180	99	18	04-.bwa.drm.sorted.bam|18	NA
chr15	20945974	40+22-	chr15	20946063	0+4-	DEL	181	99	4	04-.bwa.drm.sorted.bam|4	2608.38
chr15	20946119	40+22-	chr15	20946174	0+3-	DEL	284	99	3	04-.bwa.drm.sorted.bam|3	1547.64
chr15	21952380	26+17-	chr15	21952610	26+17-	DEL	191	99	17	04-.bwa.drm.sorted.bam|17	NA
chr15	21952610	26+17-	chr15	21952712	0+3-	DEL	210	99	3	04-.bwa.drm.sorted.bam|3	1820.75
chr15	35384540	9+5-	chr15	35384647	9+5-	ITX	-13	99	3	04-.bwa.drm.sorted.bam|3	NA
chr15	35384792	9+5-	chr15	35384853	1+3-	DEL	200	83	2	04-.bwa.drm.sorted.bam|2	8188.95
chr15	62374533	34+26-	chr15	62374731	34+26-	DEL	191	99	20	04-.bwa.drm.sorted.bam|20	NA
chr15	62374731	34+26-	chr15	62374815	0+3-	DEL	349	99	3	04-.bwa.drm.sorted.bam|3	552.73
chr15	73191496	62+32-	chr15	73191805	62+32-	DEL	206	99	29	04-.bwa.drm.sorted.bam|29	NA
chr15	73191805	62+32-	chr15	73191883	0+25-	DEL	229	99	25	04-.bwa.drm.sorted.bam|25	992.08
chr15	73191950	62+32-	chr15	73192017	0+4-	DEL	400	99	4	04-.bwa.drm.sorted.bam|4	2336.06
chr15	73454013	27+12-	chr15	73454130	27+12-	DEL	195	99	10	04-.bwa.drm.sorted.bam|10	NA
chr15	73454130	27+12-	chr15	73454194	0+15-	DEL	243	99	15	04-.bwa.drm.sorted.bam|15	2418.18
chr15	90631671	25+10-	chr15	90631981	25+10-	ITX	-12	99	5	04-.bwa.drm.sorted.bam|5	NA
chr15	92829675	29+0-	chr15	92829754	5+30-	DEL	222	99	29	04-.bwa.drm.sorted.bam|29	8619.75
chr15	92830156	31+20-	chr15	92830262	31+20-	DEL	170	99	15	04-.bwa.drm.sorted.bam|15	NA
chr15	92830262	31+20-	chr15	92830334	0+4-	DEL	250	99	4	04-.bwa.drm.sorted.bam|4	2149.50
chr16	5416426	46+36-	chr16	5416824	46+36-	DEL	222	99	36	04-.bwa.drm.sorted.bam|36	NA
chr17	7572907	21+15-	chr17	7573065	21+15-	DEL	178	99	9	04-.bwa.drm.sorted.bam|9	NA
chr17	7573947	9+0-	chr17	7574006	16+10-	DEL	179	99	6	04-.bwa.drm.sorted.bam|6	9443.21
chr17	7574176	16+10-	chr17	7574235	0+7-	DEL	200	99	7	04-.bwa.drm.sorted.bam|7	2885.43
chr17	7576245	2+0-	chr17	7576303	115+77-	DEL	205	99	67	04-.bwa.drm.sorted.bam|67	NA
chr17	7577171	115+77-	chr17	7577247	3+11-	DEL	183	99	11	04-.bwa.drm.sorted.bam|11	22400.01
chr17	7577450	12+4-	chr17	7577511	12+4-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	NA
chr17	7578201	20+6-	chr17	7578300	20+6-	DEL	173	80	2	04-.bwa.drm.sorted.bam|2	NA
chr17	7578421	19+6-	chr17	7578557	19+6-	ITX	-12	99	5	04-.bwa.drm.sorted.bam|5	NA
chr17	7578702	19+6-	chr17	7578706	0+3-	DEL	166	99	3	04-.bwa.drm.sorted.bam|3	5297.28
chr17	7579007	2+1-	chr17	7579063	34+32-	DEL	211	99	18	04-.bwa.drm.sorted.bam|18	846.97
chr17	7579007	8+0-	chr17	7579063	34+32-	DEL	257	99	8	04-.bwa.drm.sorted.bam|8	829.09
chr17	7579538	34+32-	chr17	7579613	23+16-	DEL	181	99	8	04-.bwa.drm.sorted.bam|8	11555.69
chr17	7579898	23+16-	chr17	7579953	0+2-	DEL	178	76	2	04-.bwa.drm.sorted.bam|2	8723.05
chr17	37921761	2+0-	chr17	37922269	5+5-	ITX	-13	99	3	04-.bwa.drm.sorted.bam|3	365.58
chr17	74732992	27+19-	chr17	74733232	27+19-	DEL	190	99	12	04-.bwa.drm.sorted.bam|12	NA
chr17	74733232	27+19-	chr17	74733372	0+2-	DEL	155	72	2	04-.bwa.drm.sorted.bam|2	2100.36
chr18	23785676	30+29-	chr18	23786069	30+29-	DEL	212	99	28	04-.bwa.drm.sorted.bam|28	NA
chr18	39368792	10+0-	chr18	39368850	62+66-	DEL	222	99	62	04-.bwa.drm.sorted.bam|62	266.83
chr18	42531649	6+0-	chr18	42531722	43+44-	DEL	196	99	39	04-.bwa.drm.sorted.bam|39	848.02
chr18	73424550	2+1-	chr18	73424652	0+2-	DEL	206	93	2	04-.bwa.drm.sorted.bam|2	689.23
chr19	7805315	114+102-	chr19	7805903	114+102-	DEL	218	99	91	04-.bwa.drm.sorted.bam|91	NA
chr19	7806462	34+12-	chr19	7806611	34+12-	DEL	171	99	9	04-.bwa.drm.sorted.bam|9	NA
chr19	7806611	34+12-	chr19	7806663	14+17-	DEL	195	99	15	04-.bwa.drm.sorted.bam|15	5357.21
chr19	7806868	14+17-	chr19	7806937	0+6-	DEL	221	99	6	04-.bwa.drm.sorted.bam|6	5831.68
chr19	13054281	2+0-	chr19	13054801	27+17-	ITX	-12	99	13	04-.bwa.drm.sorted.bam|13	714.29
chr19	13054656	27+17-	chr19	13054710	4+4-	DEL	168	99	4	04-.bwa.drm.sorted.bam|4	6305.19
chr19	13054943	4+4-	chr19	13054994	0+2-	DEL	183	91	2	04-.bwa.drm.sorted.bam|2	236.88
chr19	17948084	29+17-	chr19	17948312	29+17-	DEL	197	99	9	04-.bwa.drm.sorted.bam|9	NA
chr19	33792106	24+11-	chr19	33792357	24+11-	ITX	-13	99	6	04-.bwa.drm.sorted.bam|6	NA
chr19	33792357	24+11-	chr19	33792472	5+9-	DEL	195	99	8	04-.bwa.drm.sorted.bam|8	12650.25
chr19	33793070	2+1-	chr19	33793216	0+3-	DEL	189	99	2	04-.bwa.drm.sorted.bam|2	9892.11
chr19	33793027	6+4-	chr19	33793118	6+4-	ITX	-11	99	4	04-.bwa.drm.sorted.bam|4	NA
chr19	45297448	11+4-	chr19	45297621	11+4-	DEL	159	76	2	04-.bwa.drm.sorted.bam|2	NA
chr19	45297766	11+4-	chr19	45297886	0+2-	DEL	234	75	2	04-.bwa.drm.sorted.bam|2	1051.23
chr19	45303694	11+7-	chr19	45303842	11+7-	ITX	-11	99	5	04-.bwa.drm.sorted.bam|5	NA
chr20	31021851	2+0-	chr20	31021984	24+17-	DEL	177	99	15	04-.bwa.drm.sorted.bam|15	814.55
chr20	31022662	287+165-	chr20	31025266	287+165-	DEL	198	99	112	04-.bwa.drm.sorted.bam|112	NA
chr20	37606244	38+39-	chr20	37606636	38+39-	DEL	235	99	36	04-.bwa.drm.sorted.bam|36	NA
chr20	48808325	12+9-	chr20	48808569	12+9-	DEL	173	99	9	04-.bwa.drm.sorted.bam|9	NA
chr20	57484253	71+50-	chr20	57484882	71+50-	DEL	196	99	43	04-.bwa.drm.sorted.bam|43	NA
chr21	36171398	7+0-	chr21	36171469	29+14-	DEL	183	99	11	04-.bwa.drm.sorted.bam|11	4577.52
chr21	36171763	29+14-	chr21	36171894	0+6-	DEL	201	99	6	04-.bwa.drm.sorted.bam|6	1772.10
chr21	36193700	2+0-	chr21	36193757	44+37-	DEL	198	99	31	04-.bwa.drm.sorted.bam|31	1629.09
chr21	36206675	9+4-	chr21	36206788	9+4-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chr21	36231518	4+0-	chr21	36231617	18+9-	DEL	175	99	5	04-.bwa.drm.sorted.bam|5	1719.60
chr21	36231830	18+9-	chr21	36231887	22+10-	DEL	194	99	7	04-.bwa.drm.sorted.bam|7	20906.68
chr21	36231971	22+10-	chr21	36232102	0+7-	DEL	207	99	7	04-.bwa.drm.sorted.bam|7	3426.07
chr21	36232116	22+10-	chr21	36232292	0+2-	DEL	366	87	2	04-.bwa.drm.sorted.bam|2	1783.88
chr21	36252639	62+55-	chr21	36253233	62+55-	DEL	206	99	52	04-.bwa.drm.sorted.bam|52	NA
chr21	36258923	3+0-	chr21	36258996	26+17-	DEL	201	99	12	04-.bwa.drm.sorted.bam|12	4452.11
chr21	36264979	2+0-	chr21	36265043	60+58-	DEL	214	99	56	04-.bwa.drm.sorted.bam|56	483.64
chr21	36420728	2+0-	chr21	36421393	22+15-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	651.64
chr21	36420947	8+0-	chr21	36421003	22+15-	DEL	218	99	8	04-.bwa.drm.sorted.bam|8	3316.37
chr21	36421248	22+15-	chr21	36421308	0+2-	DEL	207	79	2	04-.bwa.drm.sorted.bam|2	3611.15
chr21	36421393	22+15-	chr21	36421404	0+4-	DEL	211	99	4	04-.bwa.drm.sorted.bam|4	2976.23
chr21	36971918	6+0-	chr21	36971991	44+47-	DEL	231	99	45	04-.bwa.drm.sorted.bam|45	3180.08
chr21	44514715	47+22-	chr21	44514995	47+22-	DEL	187	99	11	04-.bwa.drm.sorted.bam|11	NA
chr21	44514995	47+22-	chr21	44515061	0+12-	DEL	242	99	12	04-.bwa.drm.sorted.bam|12	1641.43
chr21	44524196	100+88-	chr21	44524574	100+88-	DEL	214	99	87	04-.bwa.drm.sorted.bam|87	NA
chr22	30290218	5+1-	chr22	30290310	0+5-	DEL	173	99	5	04-.bwa.drm.sorted.bam|5	10766.17
chr22	30293874	8+1-	chr22	30293875	0+2-	DEL	152	99	2	04-.bwa.drm.sorted.bam|2	3604.09
chr22	30293874	8+1-	chr22	30293967	0+3-	DEL	243	99	3	04-.bwa.drm.sorted.bam|3	2471.02
chrX	14852441	37+29-	chrX	14852913	37+29-	DEL	228	99	25	04-.bwa.drm.sorted.bam|25	NA
chrX	15808510	15+7-	chrX	15808710	15+7-	DEL	214	99	4	04-.bwa.drm.sorted.bam|4	NA
chrX	15808710	15+7-	chrX	15808771	11+5-	DEL	239	99	5	04-.bwa.drm.sorted.bam|5	7357.62
chrX	15808915	11+5-	chrX	15808982	30+26-	DEL	206	99	24	04-.bwa.drm.sorted.bam|24	3464.86
chrX	15809276	30+26-	chrX	15809413	0+5-	DEL	240	99	5	04-.bwa.drm.sorted.bam|5	2372.29
chrX	15817810	28+21-	chrX	15818088	28+21-	DEL	208	99	19	04-.bwa.drm.sorted.bam|19	NA
chrX	15818233	28+21-	chrX	15818297	0+2-	DEL	243	72	2	04-.bwa.drm.sorted.bam|2	1184.79
chrX	15821626	74+62-	chrX	15822571	74+62-	DEL	215	99	59	04-.bwa.drm.sorted.bam|59	NA
chrX	15826037	3+0-	chrX	15826102	45+34-	DEL	210	99	30	04-.bwa.drm.sorted.bam|30	714.29
chrX	15826682	45+34-	chrX	15826729	0+3-	DEL	255	99	3	04-.bwa.drm.sorted.bam|3	1370.30
chrX	15827159	37+21-	chrX	15827420	37+21-	DEL	201	99	19	04-.bwa.drm.sorted.bam|19	NA
chrX	15827420	37+21-	chrX	15827473	3+14-	DEL	211	99	13	04-.bwa.drm.sorted.bam|13	18396.44
chrX	15833579	6+0-	chrX	15833687	5+9-	DEL	186	99	5	04-.bwa.drm.sorted.bam|5	7164.99
chrX	15836569	31+26-	chrX	15836977	31+26-	DEL	210	99	22	04-.bwa.drm.sorted.bam|22	NA
chrX	15838114	9+0-	chrX	15838189	19+19-	DEL	239	99	15	04-.bwa.drm.sorted.bam|15	2269.87
chrX	15838458	19+19-	chrX	15838515	0+5-	DEL	184	99	5	04-.bwa.drm.sorted.bam|5	3801.21
chrX	15840617	6+0-	chrX	15840722	44+31-	DEL	219	99	28	04-.bwa.drm.sorted.bam|28	1179.15
chrX	15841423	44+31-	chrX	15841504	0+2-	DEL	252	65	2	04-.bwa.drm.sorted.bam|2	3248.13
chrX	32224685	17+15-	chrX	32224989	17+15-	DEL	201	99	14	04-.bwa.drm.sorted.bam|14	NA
chrX	32224989	17+15-	chrX	32225094	0+2-	DEL	328	71	2	04-.bwa.drm.sorted.bam|2	294.79
chrX	39911462	46+34-	chrX	39911741	46+34-	DEL	191	99	32	04-.bwa.drm.sorted.bam|32	NA
chrX	39911741	46+34-	chrX	39911810	0+4-	DEL	193	99	4	04-.bwa.drm.sorted.bam|4	224.30
chrX	39913000	8+2-	chrX	39913090	8+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	39913090	8+2-	chrX	39913153	49+31-	DEL	212	99	22	04-.bwa.drm.sorted.bam|22	4421.82
chrX	39913681	49+31-	chrX	39913741	0+7-	DEL	215	99	7	04-.bwa.drm.sorted.bam|7	2837.33
chrX	39914407	8+0-	chrX	39914483	12+12-	DEL	208	99	10	04-.bwa.drm.sorted.bam|10	2240.00
chrX	39916502	3+0-	chrX	39916581	1+3-	DEL	162	88	2	04-.bwa.drm.sorted.bam|2	4897.59
chrX	39921496	10+3-	chrX	39921632	10+3-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	NA
chrX	39921632	10+3-	chrX	39921697	2+4-	DEL	165	99	3	04-.bwa.drm.sorted.bam|3	3809.57
chrX	39921816	2+4-	chrX	39921877	19+15-	DEL	195	99	10	04-.bwa.drm.sorted.bam|10	4059.38
chrX	39922547	3+0-	chrX	39922571	11+8-	DEL	196	99	5	04-.bwa.drm.sorted.bam|5	3022.01
chrX	39922953	8+4-	chrX	39923108	8+4-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	NA
chrX	39923624	23+13-	chrX	39923938	23+13-	DEL	198	99	8	04-.bwa.drm.sorted.bam|8	NA
chrX	39930041	10+0-	chrX	39930162	106+81-	DEL	204	99	72	04-.bwa.drm.sorted.bam|72	5627.77
chrX	39931003	106+81-	chrX	39931058	4+23-	DEL	222	99	23	04-.bwa.drm.sorted.bam|23	3095.27
chrX	39931491	4+23-	chrX	39931501	48+36-	DEL	199	99	23	04-.bwa.drm.sorted.bam|23	8886.43
chrX	39931450	4+1-	chrX	39931501	48+36-	DEL	187	64	2	04-.bwa.drm.sorted.bam|2	12441.79
chrX	39932557	10+2-	chrX	39932619	10+10-	DEL	172	99	6	04-.bwa.drm.sorted.bam|6	13729.04
chrX	39932903	11+3-	chrX	39933047	11+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	39933047	11+3-	chrX	39933103	9+3-	DEL	180	99	3	04-.bwa.drm.sorted.bam|3	13541.83
chrX	39933197	9+3-	chrX	39933271	15+9-	DEL	203	99	5	04-.bwa.drm.sorted.bam|5	13803.25
chrX	39933558	15+9-	chrX	39933621	5+5-	DEL	174	99	4	04-.bwa.drm.sorted.bam|4	10317.58
chrX	39933827	4+3-	chrX	39933873	4+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	39933945	14+4-	chrX	39934097	14+4-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	39934097	14+4-	chrX	39934148	3+3-	DEL	165	81	2	04-.bwa.drm.sorted.bam|2	10621.04
chrX	39934242	14+4-	chrX	39934269	6+4-	DEL	180	77	2	04-.bwa.drm.sorted.bam|2	14396.62
chrX	39935676	23+11-	chrX	39935796	23+11-	DEL	178	99	7	04-.bwa.drm.sorted.bam|7	NA
chrX	39935796	23+11-	chrX	39935866	0+10-	DEL	222	99	9	04-.bwa.drm.sorted.bam|9	9728.00
chrX	39937213	5+3-	chrX	39937280	5+3-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	44732640	4+0-	chrX	44732745	12+8-	DEL	192	99	6	04-.bwa.drm.sorted.bam|6	6337.94
chrX	44733000	12+8-	chrX	44733144	6+7-	DEL	206	99	5	04-.bwa.drm.sorted.bam|5	7738.19
chrX	44733357	6+7-	chrX	44733514	0+2-	DEL	317	89	2	04-.bwa.drm.sorted.bam|2	1076.17
chrX	44820158	3+0-	chrX	44820291	65+58-	DEL	215	99	54	04-.bwa.drm.sorted.bam|54	232.73
chrX	44833695	3+0-	chrX	44833794	22+9-	DEL	226	99	9	04-.bwa.drm.sorted.bam|9	781.63
chrX	44834083	22+9-	chrX	44834146	0+7-	DEL	236	99	7	04-.bwa.drm.sorted.bam|7	245.66
chrX	44834228	22+9-	chrX	44834255	0+4-	DEL	341	99	4	04-.bwa.drm.sorted.bam|4	809.81
chrX	44869934	2+0-	chrX	44870023	38+43-	DEL	221	99	35	04-.bwa.drm.sorted.bam|35	925.94
chrX	44869918	6+0-	chrX	44870023	38+43-	DEL	205	99	6	04-.bwa.drm.sorted.bam|6	1179.15
chrX	44879525	6+0-	chrX	44879597	44+44-	DEL	218	99	42	04-.bwa.drm.sorted.bam|42	1504.65
chrX	44893858	10+0-	chrX	44893912	33+22-	DEL	231	99	20	04-.bwa.drm.sorted.bam|20	286.60
chrX	44894288	33+22-	chrX	44894363	4+9-	DEL	236	99	9	04-.bwa.drm.sorted.bam|9	12793.80
chrX	44896632	3+0-	chrX	44896735	34+27-	DEL	201	99	23	04-.bwa.drm.sorted.bam|23	2404.10
chrX	44897175	34+27-	chrX	44897247	0+4-	DEL	241	99	4	04-.bwa.drm.sorted.bam|4	214.95
chrX	44910905	13+0-	chrX	44910970	8+20-	DEL	186	99	12	04-.bwa.drm.sorted.bam|12	4523.86
chrX	44912743	6+0-	chrX	44912878	69+75-	DEL	219	99	70	04-.bwa.drm.sorted.bam|70	1604.96
chrX	44912826	5+0-	chrX	44912878	69+75-	DEL	212	99	5	04-.bwa.drm.sorted.bam|5	1190.49
chrX	44918045	4+0-	chrX	44918162	15+13-	DEL	205	99	9	04-.bwa.drm.sorted.bam|9	10185.30
chrX	44918457	15+13-	chrX	44918526	23+19-	DEL	222	99	18	04-.bwa.drm.sorted.bam|18	6280.27
chrX	44919072	23+19-	chrX	44919156	3+8-	DEL	316	95	3	04-.bwa.drm.sorted.bam|3	878.57
chrX	44919035	5+0-	chrX	44919156	3+8-	DEL	202	99	5	04-.bwa.drm.sorted.bam|5	1023.23
chrX	44920154	4+0-	chrX	44920287	11+4-	DEL	202	99	3	04-.bwa.drm.sorted.bam|3	465.45
chrX	44920366	11+4-	chrX	44920442	1+11-	DEL	191	99	9	04-.bwa.drm.sorted.bam|9	5294.55
chrX	44921692	86+56-	chrX	44922407	86+56-	DEL	224	99	51	04-.bwa.drm.sorted.bam|51	NA
chrX	44922407	86+56-	chrX	44922471	9+31-	DEL	220	99	27	04-.bwa.drm.sorted.bam|27	967.27
chrX	44922471	9+31-	chrX	44923072	18+5-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	1261.80
chrX	44922927	18+5-	chrX	44923001	12+4-	DEL	191	99	4	04-.bwa.drm.sorted.bam|4	8993.03
chrX	44923072	18+5-	chrX	44923220	0+8-	DEL	337	85	2	04-.bwa.drm.sorted.bam|2	12518.43
chrX	44923116	12+4-	chrX	44923220	0+8-	DEL	191	99	6	04-.bwa.drm.sorted.bam|6	4613.15
chrX	44928366	2+0-	chrX	44928462	44+35-	DEL	218	99	30	04-.bwa.drm.sorted.bam|30	483.64
chrX	44928990	44+35-	chrX	44929041	17+6-	DEL	215	99	6	04-.bwa.drm.sorted.bam|6	8496.83
chrX	44929332	17+6-	chrX	44929413	17+5-	DEL	201	99	5	04-.bwa.drm.sorted.bam|5	10508.65
chrX	44929610	17+5-	chrX	44929673	0+7-	DEL	193	99	7	04-.bwa.drm.sorted.bam|7	8352.33
chrX	44935759	33+25-	chrX	44936107	33+25-	DEL	194	99	19	04-.bwa.drm.sorted.bam|19	NA
chrX	44936107	33+25-	chrX	44936161	0+10-	DEL	238	99	10	04-.bwa.drm.sorted.bam|10	8597.98
chrX	44937338	11+0-	chrX	44937450	44+46-	DEL	224	99	45	04-.bwa.drm.sorted.bam|45	552.73
chrX	44937960	44+46-	chrX	44938012	21+13-	DEL	257	99	11	04-.bwa.drm.sorted.bam|11	297.62
chrX	44938318	21+13-	chrX	44938371	17+15-	DEL	188	99	13	04-.bwa.drm.sorted.bam|13	11680.28
chrX	44938469	17+15-	chrX	44938534	1+10-	DEL	173	99	9	04-.bwa.drm.sorted.bam|9	5952.45
chrX	44941721	38+16-	chrX	44941954	38+16-	DEL	197	99	13	04-.bwa.drm.sorted.bam|13	NA
chrX	44941954	38+16-	chrX	44942064	5+16-	DEL	246	99	16	04-.bwa.drm.sorted.bam|16	9285.82
chrX	44942179	5+16-	chrX	44942241	81+76-	DEL	247	99	73	04-.bwa.drm.sorted.bam|73	1248.09
chrX	44944972	47+33-	chrX	44945520	47+33-	DEL	234	99	32	04-.bwa.drm.sorted.bam|32	NA
chrX	44948736	3+0-	chrX	44948796	49+48-	DEL	206	99	45	04-.bwa.drm.sorted.bam|45	1031.76
chrX	44949825	5+0-	chrX	44949884	20+21-	DEL	194	99	21	04-.bwa.drm.sorted.bam|21	1049.25
chrX	44966464	3+0-	chrX	44966542	10+12-	DEL	339	99	3	04-.bwa.drm.sorted.bam|3	1318.61
chrX	44966464	8+0-	chrX	44966542	10+12-	DEL	198	99	7	04-.bwa.drm.sorted.bam|7	1388.91
chrX	44966690	10+12-	chrX	44966741	6+14-	DEL	195	99	13	04-.bwa.drm.sorted.bam|13	7283.00
chrX	44969294	17+8-	chrX	44969485	17+8-	DEL	203	99	4	04-.bwa.drm.sorted.bam|4	NA
chrX	44969485	17+8-	chrX	44969628	0+2-	DEL	182	75	2	04-.bwa.drm.sorted.bam|2	2164.53
chrX	44969630	17+8-	chrX	44969709	0+2-	DEL	219	75	2	04-.bwa.drm.sorted.bam|2	1658.18
chrX	44970571	24+13-	chrX	44970713	24+13-	DEL	182	99	12	04-.bwa.drm.sorted.bam|12	NA
chrX	44970713	24+13-	chrX	44970852	0+2-	DEL	233	76	2	04-.bwa.drm.sorted.bam|2	890.73
chrX	48649846	6+0-	chrX	48649875	0+2-	DEL	192	91	2	04-.bwa.drm.sorted.bam|2	7916.07
chrX	53423353	2+0-	chrX	53423355	9+4-	DEL	204	91	2	04-.bwa.drm.sorted.bam|2	4527.10
chrX	53426330	51+47-	chrX	53426797	51+47-	DEL	228	99	43	04-.bwa.drm.sorted.bam|43	NA
chrX	53432235	3+0-	chrX	53432322	7+5-	DEL	260	99	3	04-.bwa.drm.sorted.bam|3	2668.34
chrX	53442136	13+2-	chrX	53442202	0+4-	DEL	169	99	4	04-.bwa.drm.sorted.bam|4	4455.32
chrX	74804313	10+2-	chrX	74804413	10+2-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	74804413	10+2-	chrX	74804510	0+7-	DEL	186	99	7	04-.bwa.drm.sorted.bam|7	5265.16
chrX	76778556	21+14-	chrX	76778791	21+14-	DEL	204	99	12	04-.bwa.drm.sorted.bam|12	NA
chrX	76778791	21+14-	chrX	76778901	1+2-	DEL	170	73	2	04-.bwa.drm.sorted.bam|2	3376.66
chrX	76812525	4+0-	chrX	76812655	58+19-	DEL	243	99	16	04-.bwa.drm.sorted.bam|16	119.05
chrX	76813075	58+19-	chrX	76813138	2+34-	DEL	228	99	33	04-.bwa.drm.sorted.bam|33	14002.43
chrX	76813220	58+19-	chrX	76813453	0+4-	DEL	415	70	2	04-.bwa.drm.sorted.bam|2	8884.58
chrX	76813354	2+34-	chrX	76813453	0+4-	DEL	273	76	2	04-.bwa.drm.sorted.bam|2	468.98
chrX	76813932	2+0-	chrX	76813958	65+63-	DEL	229	99	55	04-.bwa.drm.sorted.bam|55	2081.62
chrX	76813907	4+0-	chrX	76813958	65+63-	DEL	249	99	4	04-.bwa.drm.sorted.bam|4	3338.04
chrX	76829274	4+0-	chrX	76829326	58+30-	DEL	202	99	28	04-.bwa.drm.sorted.bam|28	297.62
chrX	76829812	58+30-	chrX	76829871	23+42-	DEL	237	99	40	04-.bwa.drm.sorted.bam|40	11541.70
chrX	76845172	28+9-	chrX	76845350	28+9-	DEL	191	99	7	04-.bwa.drm.sorted.bam|7	NA
chrX	76845350	28+9-	chrX	76845406	0+20-	DEL	216	99	20	04-.bwa.drm.sorted.bam|20	3040.00
chrX	76848855	11+0-	chrX	76848906	52+50-	DEL	209	99	49	04-.bwa.drm.sorted.bam|49	1820.75
chrX	76848906	52+50-	chrX	76849636	6+5-	ITX	-12	99	3	04-.bwa.drm.sorted.bam|3	805.62
chrX	76854672	133+108-	chrX	76856163	133+108-	DEL	223	99	100	04-.bwa.drm.sorted.bam|100	NA
chrX	76856163	133+108-	chrX	76856216	0+7-	DEL	227	99	7	04-.bwa.drm.sorted.bam|7	876.02
chrX	76871926	3+0-	chrX	76871982	11+7-	DEL	239	99	5	04-.bwa.drm.sorted.bam|5	1385.94
chrX	76872250	11+7-	chrX	76872302	0+4-	DEL	166	99	3	04-.bwa.drm.sorted.bam|3	2976.23
chrX	76874033	69+67-	chrX	76874721	69+67-	DEL	216	99	63	04-.bwa.drm.sorted.bam|63	NA
chrX	76875605	2+0-	chrX	76875658	44+35-	DEL	200	99	33	04-.bwa.drm.sorted.bam|33	1168.03
chrX	76876151	44+35-	chrX	76876226	0+5-	DEL	351	99	5	04-.bwa.drm.sorted.bam|5	619.05
chrX	76888481	7+0-	chrX	76888580	53+13-	DEL	199	99	10	04-.bwa.drm.sorted.bam|10	2657.56
chrX	76888856	53+13-	chrX	76888911	36+68-	DEL	204	99	64	04-.bwa.drm.sorted.bam|64	13788.04
chrX	76889378	36+68-	chrX	76889431	0+4-	DEL	292	99	4	04-.bwa.drm.sorted.bam|4	584.01
chrX	76890084	3+0-	chrX	76890235	0+24-	DEL	297	87	2	04-.bwa.drm.sorted.bam|2	7738.19
chrX	76890169	25+3-	chrX	76890235	0+24-	DEL	175	99	23	04-.bwa.drm.sorted.bam|23	3517.36
chrX	76919964	63+57-	chrX	76920476	63+57-	DEL	232	99	56	04-.bwa.drm.sorted.bam|56	NA
chrX	76931498	2+0-	chrX	76931918	20+5-	ITX	-10	99	3	04-.bwa.drm.sorted.bam|3	110.55
chrX	76931773	20+5-	chrX	76931844	0+12-	DEL	203	99	12	04-.bwa.drm.sorted.bam|12	7411.22
chrX	76931918	20+5-	chrX	76932049	0+3-	DEL	290	99	3	04-.bwa.drm.sorted.bam|3	3869.09
chrX	76940116	14+0-	chrX	76940183	38+35-	DEL	230	99	34	04-.bwa.drm.sorted.bam|34	NA
chrX	76940665	38+35-	chrX	76940728	0+10-	DEL	260	99	10	04-.bwa.drm.sorted.bam|10	1965.25
chrX	100056189	6+1-	chrX	100056255	20+7-	DEL	202	99	6	04-.bwa.drm.sorted.bam|6	5158.79
chrX	100056458	20+7-	chrX	100056519	106+90-	DEL	213	99	79	04-.bwa.drm.sorted.bam|79	5074.22
chrX	100058142	106+90-	chrX	100058161	0+2-	DEL	252	56	2	04-.bwa.drm.sorted.bam|2	754.95
chrX	123156288	38+36-	chrX	123156713	38+36-	DEL	237	99	32	04-.bwa.drm.sorted.bam|32	NA
chrX	123159422	61+58-	chrX	123159979	61+58-	DEL	227	99	55	04-.bwa.drm.sorted.bam|55	NA
chrX	123164618	2+0-	chrX	123164679	17+9-	DEL	173	99	5	04-.bwa.drm.sorted.bam|5	1775.98
chrX	123165083	17+9-	chrX	123165120	0+2-	DEL	189	78	2	04-.bwa.drm.sorted.bam|2	1190.49
chrX	123171151	9+0-	chrX	123171202	41+38-	DEL	202	99	33	04-.bwa.drm.sorted.bam|33	2427.67
chrX	123171691	41+38-	chrX	123171823	0+2-	DEL	230	70	2	04-.bwa.drm.sorted.bam|2	1289.70
chrX	123176206	38+33-	chrX	123176646	38+33-	DEL	196	99	31	04-.bwa.drm.sorted.bam|31	NA
chrX	123178667	2+0-	chrX	123178771	44+34-	DEL	201	99	33	04-.bwa.drm.sorted.bam|33	148.81
chrX	123179408	44+34-	chrX	123179517	0+2-	DEL	292	66	2	04-.bwa.drm.sorted.bam|2	283.97
chrX	123180923	11+0-	chrX	123180983	37+45-	DEL	215	99	40	04-.bwa.drm.sorted.bam|40	515.88
chrX	123181491	37+45-	chrX	123181593	0+3-	DEL	346	96	3	04-.bwa.drm.sorted.bam|3	303.46
chrX	123182615	52+45-	chrX	123183076	52+45-	DEL	214	99	43	04-.bwa.drm.sorted.bam|43	NA
chrX	123183865	9+0-	chrX	123183924	4+6-	DEL	184	99	3	04-.bwa.drm.sorted.bam|3	5246.23
chrX	123184010	9+0-	chrX	123184018	7+8-	DEL	212	99	6	04-.bwa.drm.sorted.bam|6	10823.34
chrX	123184159	7+8-	chrX	123184277	0+2-	DEL	193	83	2	04-.bwa.drm.sorted.bam|2	2491.96
chrX	123184832	4+0-	chrX	123184898	10+17-	DEL	251	99	8	04-.bwa.drm.sorted.bam|8	3520.69
chrX	123184834	9+1-	chrX	123184898	10+17-	DEL	256	99	8	04-.bwa.drm.sorted.bam|8	3869.09
chrX	123185265	10+17-	chrX	123185390	0+3-	DEL	214	99	3	04-.bwa.drm.sorted.bam|3	495.24
chrX	123189732	38+26-	chrX	123190047	38+26-	DEL	209	99	22	04-.bwa.drm.sorted.bam|22	NA
chrX	123190047	38+26-	chrX	123190113	0+11-	DEL	207	99	11	04-.bwa.drm.sorted.bam|11	4689.81
chrX	123191536	51+17-	chrX	123191650	51+17-	DEL	175	99	12	04-.bwa.drm.sorted.bam|12	NA
chrX	123191650	51+17-	chrX	123191704	9+31-	DEL	202	99	28	04-.bwa.drm.sorted.bam|28	8884.58
chrX	123191795	51+17-	chrX	123191917	0+6-	DEL	307	75	2	04-.bwa.drm.sorted.bam|2	15070.62
chrX	123191865	9+31-	chrX	123191917	0+6-	DEL	194	99	4	04-.bwa.drm.sorted.bam|4	1488.11
chrX	123194805	6+0-	chrX	123194883	81+74-	DEL	224	99	70	04-.bwa.drm.sorted.bam|70	2976.23
chrX	123196553	17+0-	chrX	123196616	38+30-	DEL	229	99	24	04-.bwa.drm.sorted.bam|24	3439.19
chrX	123197012	38+30-	chrX	123197075	0+13-	DEL	225	99	13	04-.bwa.drm.sorted.bam|13	8106.67
chrX	123197852	5+2-	chrX	123197899	11+11-	DEL	176	99	7	04-.bwa.drm.sorted.bam|7	14589.71
chrX	123197845	8+3-	chrX	123197899	11+11-	DEL	226	99	4	04-.bwa.drm.sorted.bam|4	8311.38
chrX	123198162	11+11-	chrX	123198289	0+3-	DEL	207	99	3	04-.bwa.drm.sorted.bam|3	121.86
chrX	123199454	33+26-	chrX	123199844	33+26-	DEL	231	99	25	04-.bwa.drm.sorted.bam|25	NA
chrX	123199989	33+26-	chrX	123200026	9+4-	DEL	270	68	2	04-.bwa.drm.sorted.bam|2	2295.95
chrX	123200102	9+4-	chrX	123200209	33+25-	DEL	193	99	18	04-.bwa.drm.sorted.bam|18	5785.56
chrX	123200526	33+25-	chrX	123200591	0+4-	DEL	236	99	4	04-.bwa.drm.sorted.bam|4	2619.08
chrX	123201981	2+0-	chrX	123202071	82+76-	DEL	211	99	72	04-.bwa.drm.sorted.bam|72	171.96
chrX	123202567	82+76-	chrX	123202656	0+4-	DEL	195	99	4	04-.bwa.drm.sorted.bam|4	2260.59
chrX	123204724	5+0-	chrX	123204837	2+2-	DEL	184	90	2	04-.bwa.drm.sorted.bam|2	1232.63
chrX	123204869	5+0-	chrX	123204968	18+19-	DEL	187	99	12	04-.bwa.drm.sorted.bam|12	1966.26
chrX	123204907	2+2-	chrX	123204968	18+19-	DEL	229	73	2	04-.bwa.drm.sorted.bam|2	2537.11
chrX	123209981	27+16-	chrX	123210210	27+16-	DEL	199	99	15	04-.bwa.drm.sorted.bam|15	NA
chrX	123210210	27+16-	chrX	123210269	12+17-	DEL	240	99	14	04-.bwa.drm.sorted.bam|14	5770.85
chrX	123210519	12+17-	chrX	123210624	0+2-	DEL	320	79	2	04-.bwa.drm.sorted.bam|2	442.18
chrX	123211631	6+0-	chrX	123211695	33+34-	DEL	199	99	30	04-.bwa.drm.sorted.bam|30	3143.64
chrX	123214964	68+62-	chrX	123215582	68+62-	DEL	234	99	61	04-.bwa.drm.sorted.bam|61	NA
chrX	123215582	68+62-	chrX	123215635	0+2-	DEL	259	65	2	04-.bwa.drm.sorted.bam|2	292.01
chrX	123216933	2+0-	chrX	123217009	50+46-	DEL	237	99	43	04-.bwa.drm.sorted.bam|43	610.91
chrX	123220316	51+41-	chrX	123220801	51+41-	DEL	196	99	33	04-.bwa.drm.sorted.bam|33	NA
chrX	123224331	3+0-	chrX	123224341	52+25-	DEL	190	99	20	04-.bwa.drm.sorted.bam|20	6090.70
chrX	123224922	52+25-	chrX	123224981	2+6-	DEL	175	99	6	04-.bwa.drm.sorted.bam|6	7344.72
chrX	123224922	52+25-	chrX	123225067	0+4-	DEL	227	99	4	04-.bwa.drm.sorted.bam|4	5123.21
chrX	123227692	3+0-	chrX	123227725	31+8-	DEL	219	99	3	04-.bwa.drm.sorted.bam|3	2173.65
chrX	123227641	3+0-	chrX	123227725	31+8-	DEL	175	80	2	04-.bwa.drm.sorted.bam|2	3316.37
chrX	123227923	31+8-	chrX	123227982	3+15-	DEL	198	99	14	04-.bwa.drm.sorted.bam|14	11279.39
chrX	123229182	17+2-	chrX	123229233	10+3-	DEL	183	86	2	04-.bwa.drm.sorted.bam|2	16386.75
chrX	123229182	17+2-	chrX	123229317	9+24-	DEL	228	99	17	04-.bwa.drm.sorted.bam|17	16164.21
chrX	123229252	10+3-	chrX	123229317	9+24-	DEL	230	99	6	04-.bwa.drm.sorted.bam|6	10238.21
chrX	123234260	45+27-	chrX	123234562	45+27-	DEL	214	99	25	04-.bwa.drm.sorted.bam|25	NA
chrX	123234562	45+27-	chrX	123234648	0+15-	DEL	220	99	15	04-.bwa.drm.sorted.bam|15	1439.66
chrX	123415046	10+0-	chrX	123415109	31+38-	DEL	227	99	32	04-.bwa.drm.sorted.bam|32	1473.94
chrX	129146424	3+0-	chrX	129146429	12+9-	DEL	238	99	3	04-.bwa.drm.sorted.bam|3	3714.33
chrX	129146363	4+0-	chrX	129146429	12+9-	DEL	180	99	4	04-.bwa.drm.sorted.bam|4	6800.22
chrX	129146602	12+9-	chrX	129146657	11+7-	DEL	180	99	6	04-.bwa.drm.sorted.bam|6	5909.16
chrX	129146824	11+7-	chrX	129146879	19+13-	DEL	170	99	8	04-.bwa.drm.sorted.bam|8	14069.43
chrX	129147181	19+13-	chrX	129147241	13+8-	DEL	199	99	6	04-.bwa.drm.sorted.bam|6	18571.65
chrX	129147554	13+8-	chrX	129147690	2+3-	DEL	195	99	3	04-.bwa.drm.sorted.bam|3	15476.37
chrX	129147878	23+8-	chrX	129148274	23+8-	ITX	-12	99	4	04-.bwa.drm.sorted.bam|4	NA
chrX	129148274	23+8-	chrX	129148336	4+2-	DEL	186	73	2	04-.bwa.drm.sorted.bam|2	10234.38
chrX	129148662	11+4-	chrX	129148819	11+4-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	129148956	30+19-	chrX	129149418	30+19-	ITX	-12	99	10	04-.bwa.drm.sorted.bam|10	NA
chrX	129149492	14+3-	chrX	129149641	14+3-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	129149641	14+3-	chrX	129149716	16+16-	DEL	173	99	11	04-.bwa.drm.sorted.bam|11	5984.20
chrX	129154960	11+1-	chrX	129155018	0+3-	DEL	211	84	2	04-.bwa.drm.sorted.bam|2	8271.85
chrX	129154960	11+1-	chrX	129155093	0+5-	DEL	178	99	4	04-.bwa.drm.sorted.bam|4	5818.19
chrX	129156645	4+0-	chrX	129156768	4+4-	DEL	173	99	3	04-.bwa.drm.sorted.bam|3	5536.26
chrX	129158762	2+1-	chrX	129159224	12+10-	ITX	-11	99	5	04-.bwa.drm.sorted.bam|5	971.46
chrX	129159079	12+10-	chrX	129159154	11+6-	DEL	178	99	3	04-.bwa.drm.sorted.bam|3	13619.21
chrX	129159336	11+6-	chrX	129159400	9+9-	DEL	202	99	6	04-.bwa.drm.sorted.bam|6	10640.00
chrX	129162518	30+23-	chrX	129162751	30+23-	DEL	202	99	21	04-.bwa.drm.sorted.bam|21	NA
chrX	129162751	30+23-	chrX	129162857	7+3-	DEL	182	71	2	04-.bwa.drm.sorted.bam|2	2190.05
chrX	129162974	7+3-	chrX	129163092	0+4-	DEL	211	99	4	04-.bwa.drm.sorted.bam|4	2623.11
chrX	129171148	3+0-	chrX	129171192	12+5-	DEL	217	99	3	04-.bwa.drm.sorted.bam|3	2620.34
chrX	129171561	12+5-	chrX	129171597	0+5-	DEL	249	99	3	04-.bwa.drm.sorted.bam|3	5643.32
chrX	129171539	3+1-	chrX	129171597	0+5-	DEL	170	86	2	04-.bwa.drm.sorted.bam|2	6670.85
chrX	129172942	2+0-	chrX	129173077	0+2-	DEL	248	99	2	04-.bwa.drm.sorted.bam|2	1879.27
chrX	129172954	2+2-	chrX	129172981	2+2-	ITX	-12	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	129173166	5+2-	chrX	129173237	5+2-	ITX	-13	99	2	04-.bwa.drm.sorted.bam|2	NA
chrX	129184564	12+6-	chrX	129184739	12+6-	ITX	-11	99	3	04-.bwa.drm.sorted.bam|3	NA
chrX	129184739	12+6-	chrX	129184806	1+4-	DEL	198	99	4	04-.bwa.drm.sorted.bam|4	5312.78
chrX	129185840	18+8-	chrX	129186094	18+8-	DEL	202	99	7	04-.bwa.drm.sorted.bam|7	NA
chrX	129186094	18+8-	chrX	129186224	0+2-	DEL	201	72	2	04-.bwa.drm.sorted.bam|2	476.20
chrX	129189498	2+0-	chrX	129190243	30+18-	ITX	-12	99	10	04-.bwa.drm.sorted.bam|10	124.64
chrX	129190098	30+18-	chrX	129190153	6+10-	DEL	228	99	9	04-.bwa.drm.sorted.bam|9	10692.77
chrX	129190265	6+10-	chrX	129190405	0+4-	DEL	215	99	4	04-.bwa.drm.sorted.bam|4	2210.91
chrX	133511472	15+0-	chrX	133511536	98+97-	DEL	214	99	90	04-.bwa.drm.sorted.bam|90	7254.55
chrX	133527333	100+89-	chrX	133528173	100+89-	DEL	219	99	84	04-.bwa.drm.sorted.bam|84	NA
chrX	133547268	8+0-	chrX	133547333	85+58-	DEL	231	99	53	04-.bwa.drm.sorted.bam|53	476.20
chrX	133548021	85+58-	chrX	133548075	0+22-	DEL	262	99	22	04-.bwa.drm.sorted.bam|22	7164.99
chrX	133548919	52+52-	chrX	133549329	52+52-	DEL	223	99	47	04-.bwa.drm.sorted.bam|47	NA
chrX	133550910	2+0-	chrX	133551040	25+29-	DEL	226	99	14	04-.bwa.drm.sorted.bam|14	2251.11
chrX	133550995	2+0-	chrX	133551040	25+29-	DEL	269	71	2	04-.bwa.drm.sorted.bam|2	3095.27
chrX	133550942	8+0-	chrX	133551040	25+29-	DEL	187	99	8	04-.bwa.drm.sorted.bam|8	4579.74
chrX	133558974	4+0-	chrX	133559043	31+38-	DEL	216	99	22	04-.bwa.drm.sorted.bam|22	2169.58
chrX	133558991	10+0-	chrX	133559043	31+38-	DEL	210	99	10	04-.bwa.drm.sorted.bam|10	2678.60
chrY	9958783	3+2-	chrY	9958804	3+2-	ITX	-7	99	2	04-.bwa.drm.sorted.bam|2	NA
chrY	15409223	2+0-	chrY	15409318	23+14-	DEL	200	99	12	04-.bwa.drm.sorted.bam|12	162.91
chrY	15409586	23+14-	chrY	15409647	0+12-	DEL	208	99	12	04-.bwa.drm.sorted.bam|12	6089.06
chrY	15410958	27+0-	chrY	15411033	0+27-	DEL	202	99	27	04-.bwa.drm.sorted.bam|27	6190.55
chrY	15417174	2+0-	chrY	15417302	7+3-	DEL	286	98	2	04-.bwa.drm.sorted.bam|2	793.66
chrY	15417342	7+3-	chrY	15417393	1+10-	DEL	203	99	5	04-.bwa.drm.sorted.bam|5	3641.50
chrY	15417369	5+0-	chrY	15417393	1+10-	DEL	235	99	5	04-.bwa.drm.sorted.bam|5	6227.18
chrY	15435261	7+0-	chrY	15435330	28+31-	DEL	208	99	27	04-.bwa.drm.sorted.bam|27	1345.77
chrY	15435671	28+31-	chrY	15435731	0+3-	DEL	227	99	3	04-.bwa.drm.sorted.bam|3	773.82
chrY	15436422	28+16-	chrY	15436617	28+16-	DEL	195	99	16	04-.bwa.drm.sorted.bam|16	NA
chrY	15436617	28+16-	chrY	15436715	0+7-	DEL	222	99	7	04-.bwa.drm.sorted.bam|7	3000.52
chrY	15436762	28+16-	chrY	15436818	0+2-	DEL	293	74	2	04-.bwa.drm.sorted.bam|2	1924.92
chrY	15437902	3+0-	chrY	15437989	15+6-	DEL	186	99	6	04-.bwa.drm.sorted.bam|6	533.67
chrY	15438211	15+6-	chrY	15438282	0+9-	DEL	180	99	9	04-.bwa.drm.sorted.bam|9	1525.84
chrY	15447738	8+4-	chrY	15447815	8+4-	DEL	169	99	3	04-.bwa.drm.sorted.bam|3	NA
chrY	15471595	2+0-	chrY	15471673	3+6-	DEL	251	82	2	04-.bwa.drm.sorted.bam|2	1179.81
chrY	15478250	3+2-	chrY	15478314	0+3-	DEL	178	89	2	04-.bwa.drm.sorted.bam|2	1426.90
chrY	15522812	17+2-	chrY	15522920	17+2-	ITX	-11	99	2	04-.bwa.drm.sorted.bam|2	NA
chrY	15522997	17+2-	chrY	15523006	0+6-	DEL	185	99	6	04-.bwa.drm.sorted.bam|6	5578.69
chrY	15522997	17+2-	chrY	15523114	0+4-	DEL	242	99	4	04-.bwa.drm.sorted.bam|4	3270.78
chrY	15581791	32+31-	chrY	15582228	32+31-	DEL	214	99	29	04-.bwa.drm.sorted.bam|29	NA
chrY	21636034	2+0-	chrY	21636143	0+3-	DEL	204	95	2	04-.bwa.drm.sorted.bam|2	5907.65
chrY	21645365	3+0-	chrY	21645460	5+8-	DEL	257	99	4	04-.bwa.drm.sorted.bam|4	2789.35
chrY	21645389	3+0-	chrY	21645460	5+8-	DEL	175	99	3	04-.bwa.drm.sorted.bam|3	5885.38
chrUn_gl000232	5011	2+0-	chrUn_gl000232	5084	18+14-	DEL	215	99	14	04-.bwa.drm.sorted.bam|14	212.01
